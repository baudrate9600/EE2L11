configuration sqi_controller_synthesised_cfg of sqi_controller is
   for synthesised
   end for;
end sqi_controller_synthesised_cfg;
