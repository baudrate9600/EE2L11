library IEEE;
use IEEE.std_logic_1164.ALL;

entity memory_tb is
end memory_tb;

