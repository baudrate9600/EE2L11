configuration counter16_behaviour_cfg of counter16 is
   for behaviour
   end for;
end counter16_behaviour_cfg;
