configuration sqi_controller_behaviour_cfg of sqi_controller is
   for behaviour
   end for;
end sqi_controller_behaviour_cfg;
