library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of sqi is
	type sqi_statae is (START, SENDING, READING, DONE);
begin
	process (clk) 
	begin

	end process;
end behaviour;

