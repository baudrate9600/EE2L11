
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture routed of memory is

  component DEL01BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL1BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD5BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component CKND2BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component CKBD12BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD8BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component LHQD1BWP7T
    port(D, E : in std_logic; Q : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component AOI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AOI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component OAI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component INVD5BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component AO221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component AOI33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component LHD1BWP7T
    port(D, E : in std_logic; Q, QN : out std_logic);
  end component;

  component OA21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component LND1BWP7T
    port(D, EN : in std_logic; Q, QN : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AO222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; Z : out std_logic);
  end component;

  component AOI211XD0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IOA21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component ND4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component OA22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component OA221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component IND3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AOI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component OA211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component MOAI22D1BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component LNQD1BWP7T
    port(D, EN : in std_logic; Q : out std_logic);
  end component;

  component OR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component IOA21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component ND2D5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component INR3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CN, CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component DFKCNQD1BWP7T
    port(CN, CP, D : in std_logic; Q : out std_logic);
  end component;

  component CKND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component DFD1BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component DFKCND0BWP7T
    port(CN, CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component TIELBWP7T
    port(ZN : out std_logic);
  end component;

  signal FE_PHN199_framebuffer_buf_150_3045, FE_PHN198_framebuffer_buf_101_2996, FE_PHN197_framebuffer_buf_106_3001, FE_PHN196_framebuffer_buf_79_2974, FE_PHN195_framebuffer_buf_126_3021 : std_logic;
  signal FE_PHN194_framebuffer_buf_118_3013, FE_PHN193_framebuffer_buf_80_2975, FE_PHN192_framebuffer_buf_133_3028, FE_PHN191_framebuffer_buf_128_3023, FE_PHN190_framebuffer_buf_154_3049 : std_logic;
  signal FE_PHN189_framebuffer_buf_155_3050, FE_PHN188_calc_buf_out_2_2873, FE_PHN187_framebuffer_buf_93_2988, FE_PHN186_calc_buf_out_8_2879, FE_PHN185_framebuffer_buf_24_2919 : std_logic;
  signal FE_PHN184_framebuffer_buf_106_3001, FE_PHN183_framebuffer_buf_101_2996, FE_PHN182_framebuffer_buf_131_3026, FE_PHN181_framebuffer_buf_104_2999, FE_PHN180_framebuffer_buf_119_3014 : std_logic;
  signal FE_PHN179_framebuffer_buf_89_2984, FE_PHN178_framebuffer_buf_4_2899, FE_PHN177_framebuffer_buf_155_3050, FE_PHN176_calc_buf_out_8_2879, FE_PHN175_framebuffer_buf_133_3028 : std_logic;
  signal FE_PHN174_framebuffer_buf_80_2975, FE_PHN173_framebuffer_buf_127_3022, FE_PHN172_framebuffer_buf_128_3023, FE_PHN171_framebuffer_buf_150_3045, FE_PHN170_framebuffer_buf_126_3021 : std_logic;
  signal FE_PHN169_framebuffer_buf_71_2966, FE_PHN168_framebuffer_buf_146_3041, FE_PHN167_framebuffer_buf_93_2988, FE_PHN166_framebuffer_buf_5_2900, FE_PHN165_framebuffer_buf_152_3047 : std_logic;
  signal FE_PHN164_calc_buf_out_13_2884, FE_PHN163_framebuffer_buf_84_2979, FE_PHN162_calc_buf_out_2_2873, FE_PHN161_framebuffer_buf_99_2994, FE_PHN160_framebuffer_buf_40_2935 : std_logic;
  signal FE_PHN159_framebuffer_buf_122_3017, FE_PHN158_framebuffer_buf_86_2981, FE_PHN157_framebuffer_buf_79_2974, FE_PHN156_framebuffer_buf_103_2998, FE_PHN155_framebuffer_buf_154_3049 : std_logic;
  signal FE_PHN154_framebuffer_buf_70_2965, FE_PHN153_framebuffer_buf_53_2948, FE_PHN152_calc_buf_out_21_2892, FE_PHN151_framebuffer_buf_120_3015, FE_PHN150_framebuffer_buf_118_3013 : std_logic;
  signal FE_PHN149_framebuffer_buf_49_2944, FE_PHN148_framebuffer_buf_157_3052, FE_PHN147_framebuffer_buf_156_3051, FE_PHN146_framebuffer_buf_55_2950, FE_PHN145_framebuffer_buf_47_2942 : std_logic;
  signal FE_PHN144_framebuffer_buf_44_2939, FE_PHN143_framebuffer_buf_37_2932, FE_PHN142_framebuffer_buf_78_2973, FE_PHN141_framebuffer_buf_132_3027, FE_PHN140_framebuffer_buf_43_2938 : std_logic;
  signal FE_PHN139_framebuffer_buf_143_3038, FE_PHN138_framebuffer_buf_88_2983, FE_PHN137_framebuffer_buf_129_3024, FE_PHN136_framebuffer_buf_12_2907, FE_PHN135_calc_buf_out_18_2889 : std_logic;
  signal FE_PHN134_framebuffer_buf_13_2908, FE_PHN133_framebuffer_buf_14_2909, FE_PHN132_framebuffer_buf_124_3019, FE_PHN131_framebuffer_buf_72_2967, FE_PHN130_framebuffer_buf_83_2978 : std_logic;
  signal FE_PHN129_framebuffer_buf_96_2991, FE_PHN128_framebuffer_buf_62_2957, FE_PHN127_framebuffer_buf_142_3037, FE_PHN126_framebuffer_buf_153_3048, FE_PHN125_framebuffer_buf_149_3044 : std_logic;
  signal FE_PHN124_framebuffer_buf_76_2971, FE_PHN123_framebuffer_buf_111_3006, FE_PHN122_framebuffer_buf_112_3007, FE_PHN121_framebuffer_buf_134_3029, FE_PHN120_framebuffer_buf_147_3042 : std_logic;
  signal FE_PHN119_framebuffer_buf_130_3025, FE_PHN118_framebuffer_buf_114_3009, FE_PHN117_framebuffer_buf_27_2922, FE_PHN116_framebuffer_buf_144_3039, FE_PHN115_framebuffer_buf_105_3000 : std_logic;
  signal FE_PHN114_framebuffer_buf_113_3008, FE_PHN113_framebuffer_buf_98_2993, FE_PHN112_framebuffer_buf_33_2928, FE_PHN111_framebuffer_buf_6_2901, FE_PHN110_framebuffer_buf_87_2982 : std_logic;
  signal FE_PHN109_framebuffer_buf_17_2912, FE_PHN108_framebuffer_buf_63_2958, FE_PHN107_framebuffer_buf_67_2962, FE_PHN106_framebuffer_buf_46_2941, FE_PHN105_framebuffer_buf_77_2972 : std_logic;
  signal FE_PHN104_framebuffer_buf_65_2960, FE_PHN103_framebuffer_buf_110_3005, FE_PHN102_framebuffer_buf_141_3036, FE_PHN101_framebuffer_buf_8_2903, FE_PHN100_framebuffer_buf_42_2937 : std_logic;
  signal FE_PHN99_framebuffer_buf_52_2947, FE_PHN98_framebuffer_buf_15_2910, FE_PHN97_framebuffer_buf_137_3032, FE_PHN96_framebuffer_buf_39_2934, FE_PHN95_framebuffer_buf_19_2914 : std_logic;
  signal FE_PHN94_calc_buf_out_19_2890, FE_PHN93_framebuffer_buf_75_2970, FE_PHN92_framebuffer_buf_145_3040, FE_PHN91_framebuffer_buf_51_2946, FE_PHN90_framebuffer_buf_34_2929 : std_logic;
  signal FE_PHN89_framebuffer_buf_69_2964, FE_PHN88_framebuffer_buf_48_2943, FE_PHN87_framebuffer_buf_58_2953, FE_PHN86_framebuffer_buf_25_2920, FE_PHN85_framebuffer_buf_16_2911 : std_logic;
  signal FE_PHN84_calc_buf_out_7_2878, FE_PHN83_calc_buf_out_6_2877, FE_PHN82_framebuffer_buf_18_2913, FE_PHN81_framebuffer_buf_140_3035, FE_PHN80_framebuffer_buf_64_2959 : std_logic;
  signal FE_PHN79_framebuffer_buf_95_2990, FE_PHN78_framebuffer_buf_109_3004, FE_PHN77_framebuffer_buf_148_3043, FE_PHN76_framebuffer_buf_22_2917, FE_PHN75_calc_buf_out_14_2885 : std_logic;
  signal FE_PHN74_framebuffer_buf_68_2963, FE_PHN73_framebuffer_buf_151_3046, FE_PHN72_framebuffer_buf_60_2955, FE_PHN71_framebuffer_buf_136_3031, FE_PHN70_framebuffer_buf_36_2931 : std_logic;
  signal FE_PHN69_framebuffer_buf_28_2923, FE_PHN68_calc_buf_out_10_2881, FE_PHN67_framebuffer_buf_21_2916, FE_PHN66_framebuffer_buf_41_2936, FE_PHN65_framebuffer_buf_56_2951 : std_logic;
  signal FE_PHN64_calc_buf_out_15_2886, FE_PHN63_framebuffer_buf_73_2968, FE_PHN62_framebuffer_buf_123_3018, FE_PHN61_framebuffer_buf_108_3003, FE_PHN60_framebuffer_buf_102_2997 : std_logic;
  signal FE_PHN59_framebuffer_buf_139_3034, FE_PHN58_framebuffer_buf_94_2989, FE_PHN57_framebuffer_buf_35_2930, FE_PHN56_framebuffer_buf_138_3033, FE_PHN55_framebuffer_buf_97_2992 : std_logic;
  signal FE_PHN54_framebuffer_buf_115_3010, FE_PHN53_framebuffer_buf_11_2906, FE_PHN52_framebuffer_buf_45_2940, FE_PHN51_framebuffer_buf_50_2945, FE_PHN50_framebuffer_buf_135_3030 : std_logic;
  signal FE_PHN49_calc_buf_out_11_2882, FE_PHN48_framebuffer_buf_66_2961, FE_PHN47_framebuffer_buf_74_2969, FE_PHN46_framebuffer_buf_125_3020, FE_PHN45_framebuffer_buf_9_2904 : std_logic;
  signal FE_PHN44_framebuffer_buf_31_2926, FE_PHN43_framebuffer_buf_1_2896, FE_PHN42_framebuffer_buf_107_3002, FE_PHN41_framebuffer_buf_26_2921, FE_PHN40_framebuffer_buf_0_2895 : std_logic;
  signal FE_PHN39_framebuffer_buf_54_2949, FE_PHN38_framebuffer_buf_10_2905, FE_PHN37_calc_buf_out_5_2876, FE_PHN36_framebuffer_buf_23_2918, FE_PHN35_framebuffer_buf_38_2933 : std_logic;
  signal FE_PHN34_framebuffer_buf_32_2927, FE_PHN33_framebuffer_buf_121_3016, FE_PHN32_calc_buf_out_12_2883, FE_PHN31_calc_buf_out_22_2893, FE_PHN30_calc_buf_out_4_2875 : std_logic;
  signal FE_PHN29_framebuffer_buf_92_2987, FE_PHN28_calc_buf_out_3_2874, FE_PHN27_framebuffer_buf_57_2952, FE_PHN26_framebuffer_buf_100_2995, FE_PHN25_calc_buf_out_20_2891 : std_logic;
  signal FE_PHN24_framebuffer_buf_61_2956, FE_PHN23_calc_buf_out_23_2894, FE_PHN22_framebuffer_buf_30_2925, FE_PHN21_framebuffer_buf_2_2897, FE_PHN20_framebuffer_buf_29_2924 : std_logic;
  signal FE_PHN19_framebuffer_buf_3_2898, FE_PHN18_framebuffer_buf_20_2915, FE_PHN17_calc_buf_out_17_2888, FE_PHN16_calc_buf_out_9_2880, FE_PHN15_calc_buf_out_16_2887 : std_logic;
  signal FE_PHN14_calc_buf_out_1_2872, FE_PHN13_calc_buf_out_0_2871, FE_PHN12_framebuffer_buf_90_2985, FE_PHN11_framebuffer_buf_91_2986, FE_PHN10_framebuffer_buf_82_2977 : std_logic;
  signal FE_PHN9_framebuffer_buf_7_2902, FE_PHN8_framebuffer_buf_85_2980, FE_PHN7_framebuffer_buf_81_2976, FE_PHN6_framebuffer_buf_59_2954, FE_RN_1 : std_logic;
  signal FE_OFN4_framebuffer_buf_116, FE_OFN3_n_0, FE_OFN2_n_0, FE_OFN1_n_0, FE_OFN0_n_0 : std_logic;
  signal CTS_16, CTS_15, CTS_14, CTS_13 : std_logic;
  signal new_sqi_address : std_logic_vector(14 downto 0);
  signal counter : std_logic_vector(7 downto 0);
  signal new_counter : std_logic_vector(7 downto 0);
  signal row_buf : std_logic_vector(5 downto 0);
  signal state : std_logic_vector(3 downto 0);
  signal new_row_buf : std_logic_vector(5 downto 0);
  signal UNCONNECTED, UNCONNECTED0, UNCONNECTED1, UNCONNECTED2, UNCONNECTED3 : std_logic;
  signal UNCONNECTED4, UNCONNECTED5, UNCONNECTED6, UNCONNECTED7, UNCONNECTED8 : std_logic;
  signal UNCONNECTED9, UNCONNECTED10, UNCONNECTED11, UNCONNECTED12, UNCONNECTED13 : std_logic;
  signal UNCONNECTED14, UNCONNECTED15, UNCONNECTED16, UNCONNECTED17, UNCONNECTED18 : std_logic;
  signal UNCONNECTED19, UNCONNECTED20, UNCONNECTED21, UNCONNECTED22, UNCONNECTED23 : std_logic;
  signal calc_buf_out_0_2871, calc_buf_out_1_2872, calc_buf_out_2_2873, calc_buf_out_3_2874, calc_buf_out_4_2875 : std_logic;
  signal calc_buf_out_5_2876, calc_buf_out_6_2877, calc_buf_out_7_2878, calc_buf_out_8_2879, calc_buf_out_9_2880 : std_logic;
  signal calc_buf_out_10_2881, calc_buf_out_11_2882, calc_buf_out_12_2883, calc_buf_out_13_2884, calc_buf_out_14_2885 : std_logic;
  signal calc_buf_out_15_2886, calc_buf_out_16_2887, calc_buf_out_17_2888, calc_buf_out_18_2889, calc_buf_out_19_2890 : std_logic;
  signal calc_buf_out_20_2891, calc_buf_out_21_2892, calc_buf_out_22_2893, calc_buf_out_23_2894, framebuffer_buf_0_2895 : std_logic;
  signal framebuffer_buf_1_2896, framebuffer_buf_2_2897, framebuffer_buf_3_2898, framebuffer_buf_4_2899, framebuffer_buf_5_2900 : std_logic;
  signal framebuffer_buf_6_2901, framebuffer_buf_7_2902, framebuffer_buf_8_2903, framebuffer_buf_9_2904, framebuffer_buf_10_2905 : std_logic;
  signal framebuffer_buf_11_2906, framebuffer_buf_12_2907, framebuffer_buf_13_2908, framebuffer_buf_14_2909, framebuffer_buf_15_2910 : std_logic;
  signal framebuffer_buf_16_2911, framebuffer_buf_17_2912, framebuffer_buf_18_2913, framebuffer_buf_19_2914, framebuffer_buf_20_2915 : std_logic;
  signal framebuffer_buf_21_2916, framebuffer_buf_22_2917, framebuffer_buf_23_2918, framebuffer_buf_24_2919, framebuffer_buf_25_2920 : std_logic;
  signal framebuffer_buf_26_2921, framebuffer_buf_27_2922, framebuffer_buf_28_2923, framebuffer_buf_29_2924, framebuffer_buf_30_2925 : std_logic;
  signal framebuffer_buf_31_2926, framebuffer_buf_32_2927, framebuffer_buf_33_2928, framebuffer_buf_34_2929, framebuffer_buf_35_2930 : std_logic;
  signal framebuffer_buf_36_2931, framebuffer_buf_37_2932, framebuffer_buf_38_2933, framebuffer_buf_39_2934, framebuffer_buf_40_2935 : std_logic;
  signal framebuffer_buf_41_2936, framebuffer_buf_42_2937, framebuffer_buf_43_2938, framebuffer_buf_44_2939, framebuffer_buf_45_2940 : std_logic;
  signal framebuffer_buf_46_2941, framebuffer_buf_47_2942, framebuffer_buf_48_2943, framebuffer_buf_49_2944, framebuffer_buf_50_2945 : std_logic;
  signal framebuffer_buf_51_2946, framebuffer_buf_52_2947, framebuffer_buf_53_2948, framebuffer_buf_54_2949, framebuffer_buf_55_2950 : std_logic;
  signal framebuffer_buf_56_2951, framebuffer_buf_57_2952, framebuffer_buf_58_2953, framebuffer_buf_59_2954, framebuffer_buf_60_2955 : std_logic;
  signal framebuffer_buf_61_2956, framebuffer_buf_62_2957, framebuffer_buf_63_2958, framebuffer_buf_64_2959, framebuffer_buf_65_2960 : std_logic;
  signal framebuffer_buf_66_2961, framebuffer_buf_67_2962, framebuffer_buf_68_2963, framebuffer_buf_69_2964, framebuffer_buf_70_2965 : std_logic;
  signal framebuffer_buf_71_2966, framebuffer_buf_72_2967, framebuffer_buf_73_2968, framebuffer_buf_74_2969, framebuffer_buf_75_2970 : std_logic;
  signal framebuffer_buf_76_2971, framebuffer_buf_77_2972, framebuffer_buf_78_2973, framebuffer_buf_79_2974, framebuffer_buf_80_2975 : std_logic;
  signal framebuffer_buf_81_2976, framebuffer_buf_82_2977, framebuffer_buf_83_2978, framebuffer_buf_84_2979, framebuffer_buf_85_2980 : std_logic;
  signal framebuffer_buf_86_2981, framebuffer_buf_87_2982, framebuffer_buf_88_2983, framebuffer_buf_89_2984, framebuffer_buf_90_2985 : std_logic;
  signal framebuffer_buf_91_2986, framebuffer_buf_92_2987, framebuffer_buf_93_2988, framebuffer_buf_94_2989, framebuffer_buf_95_2990 : std_logic;
  signal framebuffer_buf_96_2991, framebuffer_buf_97_2992, framebuffer_buf_98_2993, framebuffer_buf_99_2994, framebuffer_buf_100_2995 : std_logic;
  signal framebuffer_buf_101_2996, framebuffer_buf_102_2997, framebuffer_buf_103_2998, framebuffer_buf_104_2999, framebuffer_buf_105_3000 : std_logic;
  signal framebuffer_buf_106_3001, framebuffer_buf_107_3002, framebuffer_buf_108_3003, framebuffer_buf_109_3004, framebuffer_buf_110_3005 : std_logic;
  signal framebuffer_buf_111_3006, framebuffer_buf_112_3007, framebuffer_buf_113_3008, framebuffer_buf_114_3009, framebuffer_buf_115_3010 : std_logic;
  signal framebuffer_buf_118_3013, framebuffer_buf_119_3014, framebuffer_buf_120_3015, framebuffer_buf_121_3016, framebuffer_buf_122_3017 : std_logic;
  signal framebuffer_buf_123_3018, framebuffer_buf_124_3019, framebuffer_buf_125_3020, framebuffer_buf_126_3021, framebuffer_buf_127_3022 : std_logic;
  signal framebuffer_buf_128_3023, framebuffer_buf_129_3024, framebuffer_buf_130_3025, framebuffer_buf_131_3026, framebuffer_buf_132_3027 : std_logic;
  signal framebuffer_buf_133_3028, framebuffer_buf_134_3029, framebuffer_buf_135_3030, framebuffer_buf_136_3031, framebuffer_buf_137_3032 : std_logic;
  signal framebuffer_buf_138_3033, framebuffer_buf_139_3034, framebuffer_buf_140_3035, framebuffer_buf_141_3036, framebuffer_buf_142_3037 : std_logic;
  signal framebuffer_buf_143_3038, framebuffer_buf_144_3039, framebuffer_buf_145_3040, framebuffer_buf_146_3041, framebuffer_buf_147_3042 : std_logic;
  signal framebuffer_buf_148_3043, framebuffer_buf_149_3044, framebuffer_buf_150_3045, framebuffer_buf_151_3046, framebuffer_buf_152_3047 : std_logic;
  signal framebuffer_buf_153_3048, framebuffer_buf_154_3049, framebuffer_buf_155_3050, framebuffer_buf_156_3051, framebuffer_buf_157_3052 : std_logic;
  signal n_0, n_1, n_2, n_3, n_4 : std_logic;
  signal n_5, n_6, n_7, n_8, n_9 : std_logic;
  signal n_10, n_11, n_12, n_13, n_14 : std_logic;
  signal n_15, n_16, n_17, n_18, n_19 : std_logic;
  signal n_20, n_21, n_22, n_23, n_24 : std_logic;
  signal n_25, n_26, n_27, n_28, n_29 : std_logic;
  signal n_30, n_31, n_32, n_33, n_34 : std_logic;
  signal n_35, n_36, n_37, n_38, n_39 : std_logic;
  signal n_40, n_41, n_42, n_43, n_44 : std_logic;
  signal n_45, n_46, n_47, n_48, n_49 : std_logic;
  signal n_50, n_51, n_53, n_54, n_55 : std_logic;
  signal n_56, n_57, n_58, n_59, n_60 : std_logic;
  signal n_61, n_62, n_63, n_64, n_65 : std_logic;
  signal n_66, n_67, n_68, n_69, n_70 : std_logic;
  signal n_71, n_72, n_73, n_74, n_75 : std_logic;
  signal n_76, n_77, n_78, n_79, n_80 : std_logic;
  signal n_81, n_82, n_83, n_84, n_85 : std_logic;
  signal n_86, n_87, n_88, n_89, n_90 : std_logic;
  signal n_91, n_92, n_93, n_95, n_97 : std_logic;
  signal n_99, n_100, n_101, n_102, n_103 : std_logic;
  signal n_105, n_106, n_107, n_108, n_109 : std_logic;
  signal n_110, n_111, n_112, n_113, n_114 : std_logic;
  signal n_115, n_116, n_117, n_118, n_119 : std_logic;
  signal n_120, n_121, n_122, n_123, n_124 : std_logic;
  signal n_125, n_126, n_127, n_128, n_129 : std_logic;
  signal n_130, n_131, n_132, n_133, n_134 : std_logic;
  signal n_135, n_136, n_137, n_138, n_139 : std_logic;
  signal n_140, n_141, n_142, n_143, n_144 : std_logic;
  signal n_145, n_146, n_147, n_148, n_150 : std_logic;
  signal n_151, n_152, n_153, n_155, n_156 : std_logic;
  signal n_157, n_158, n_159, n_160, n_161 : std_logic;
  signal n_162, n_163, n_164, n_165, n_166 : std_logic;
  signal n_167, n_168, n_169, n_170, n_171 : std_logic;
  signal n_172, n_173, n_174, n_175, n_176 : std_logic;
  signal n_177, n_178, n_179, n_180, n_181 : std_logic;
  signal n_182, n_183, n_184, n_185, n_186 : std_logic;
  signal n_187, n_188, n_189, n_190, n_191 : std_logic;
  signal n_192, n_193, n_194, n_195, n_196 : std_logic;
  signal n_197, n_198, n_199, n_200, n_202 : std_logic;
  signal n_203, n_204, n_205, n_206, n_207 : std_logic;
  signal n_208, n_209, n_210, n_211, n_212 : std_logic;
  signal n_213, n_214, n_215, n_216, n_217 : std_logic;
  signal n_218, n_219, n_221, n_222, n_223 : std_logic;
  signal n_224, n_225, n_226, n_227, n_228 : std_logic;
  signal n_229, n_230, n_231, n_232, n_233 : std_logic;
  signal n_234, n_235, n_236, n_237, n_238 : std_logic;
  signal n_239, n_240, n_241, n_242, n_243 : std_logic;
  signal n_244, n_245, n_246, n_247, n_248 : std_logic;
  signal n_250, n_251, n_252, n_253, n_254 : std_logic;
  signal n_255, n_256, n_257, n_258, n_259 : std_logic;
  signal n_261, n_262, n_263, n_264, n_265 : std_logic;
  signal n_267, n_268, n_269, n_270, n_271 : std_logic;
  signal n_272, n_273, n_274, n_275, n_276 : std_logic;
  signal n_277, n_278, n_279, n_280, n_281 : std_logic;
  signal n_283, n_284, n_285, n_286, n_287 : std_logic;
  signal n_289, n_290, n_291, n_292, n_293 : std_logic;
  signal n_294, n_295, n_296, n_297, n_298 : std_logic;
  signal n_299, n_301, n_302, n_303, n_305 : std_logic;
  signal n_306, n_307, n_308, n_309, n_310 : std_logic;
  signal n_311, n_312, n_313, n_314, n_315 : std_logic;
  signal n_316, n_317, n_318, n_319, n_320 : std_logic;
  signal n_321, n_323, n_324, n_325, n_326 : std_logic;
  signal n_327, n_328, n_329, n_330, n_331 : std_logic;
  signal n_332, n_333, n_334, n_335, n_336 : std_logic;
  signal n_337, n_338, n_339, n_340, n_341 : std_logic;
  signal n_342, n_343, n_344, n_345, n_346 : std_logic;
  signal n_347, n_348, n_350, n_351, n_352 : std_logic;
  signal n_353, n_354, n_355, n_356, n_357 : std_logic;
  signal n_358, n_359, n_360, n_361, n_362 : std_logic;
  signal n_363, n_364, n_365, n_366, n_367 : std_logic;
  signal n_368, n_369, n_370, n_371, n_372 : std_logic;
  signal n_373, n_374, n_375, n_376, n_377 : std_logic;
  signal n_378, n_379, n_380, n_381, n_382 : std_logic;
  signal n_383, n_384, n_385, n_386, n_387 : std_logic;
  signal n_388, n_389, n_390, n_391, n_392 : std_logic;
  signal n_393, n_396, n_397, n_398, n_399 : std_logic;
  signal n_400, n_401, n_402, n_403, n_404 : std_logic;
  signal n_405, n_406, n_408, n_409, n_410 : std_logic;
  signal n_411, n_418, n_419, n_420, n_421 : std_logic;
  signal n_422, n_423, n_424, n_425, n_426 : std_logic;
  signal n_427, n_428, n_429, n_430, n_431 : std_logic;
  signal n_432, n_433, n_434, n_435, n_436 : std_logic;
  signal n_437, n_438, n_439, n_440, n_441 : std_logic;
  signal n_442, n_443, n_444, n_445, n_446 : std_logic;
  signal n_447, n_448, n_449, n_450, n_451 : std_logic;
  signal n_452, n_453, n_454, n_455, n_456 : std_logic;
  signal n_457, n_459, n_460, n_461, n_462 : std_logic;
  signal n_463, n_464, n_465, n_466, n_467 : std_logic;
  signal n_468, n_469, n_470, n_471, n_472 : std_logic;
  signal n_473, n_474, n_475, n_476, n_477 : std_logic;
  signal n_478, n_479, n_483, n_484, n_485 : std_logic;
  signal n_486, n_488, n_489, n_490, n_491 : std_logic;
  signal n_492, n_493, n_494, n_495, n_496 : std_logic;
  signal n_497, n_498, n_499, n_500, n_501 : std_logic;
  signal n_502, n_503, n_504, n_505, n_506 : std_logic;
  signal n_507, n_508, n_509, n_510, n_511 : std_logic;
  signal n_512, n_513, n_514, n_515, n_516 : std_logic;
  signal n_517, n_518, n_519, n_520, n_521 : std_logic;
  signal n_522, n_523, n_524, n_525, n_526 : std_logic;
  signal n_527, n_528, n_529, n_530, n_531 : std_logic;
  signal n_532, n_533, n_534, n_535, n_536 : std_logic;
  signal n_537, n_538, n_539, n_540, n_541 : std_logic;
  signal n_542, n_543, n_544, n_545, n_546 : std_logic;
  signal n_547, n_548, n_549, n_550, n_551 : std_logic;
  signal n_552, n_553, n_554, n_555, n_556 : std_logic;
  signal n_557, n_558, n_559, n_560, n_561 : std_logic;
  signal n_562, n_563, n_564, n_565, n_566 : std_logic;
  signal n_567, n_568, n_569, n_570, n_571 : std_logic;
  signal n_572, n_573, n_574, n_575, n_576 : std_logic;
  signal n_577, n_578, n_579, n_580, n_581 : std_logic;
  signal n_582, n_583, n_584, n_585, n_586 : std_logic;
  signal n_587, n_588, n_589, n_590, n_591 : std_logic;
  signal n_592, n_593, n_594, n_595, n_596 : std_logic;
  signal n_597, n_598, n_599, n_600, n_601 : std_logic;
  signal n_602, n_603, n_604, n_605, n_606 : std_logic;
  signal n_607, n_608, n_609, n_610, n_611 : std_logic;
  signal n_612, n_613, n_614, n_615, n_616 : std_logic;
  signal n_617, n_618, n_619, n_620, n_621 : std_logic;
  signal n_622, n_623, n_624, n_625, n_626 : std_logic;
  signal n_627, n_628, n_629, n_630, n_631 : std_logic;
  signal n_632, n_633, n_634, n_635, n_636 : std_logic;
  signal n_637, n_638, n_639, n_640, n_641 : std_logic;
  signal n_642, n_643, n_644, n_645, n_646 : std_logic;
  signal n_647, n_648, n_649, n_650, n_651 : std_logic;
  signal n_652, n_653, n_654, n_655, n_656 : std_logic;
  signal n_657, n_658, n_659, n_660, n_661 : std_logic;
  signal n_662, n_664, n_665, n_666, n_667 : std_logic;
  signal n_668, n_669, n_670, n_671, n_672 : std_logic;
  signal n_674, n_675, n_676, n_677, n_678 : std_logic;
  signal n_679, n_680, n_681, n_682, n_684 : std_logic;
  signal n_685, n_686, n_687, n_688, n_689 : std_logic;
  signal n_690, n_691, n_692, n_693, n_694 : std_logic;
  signal n_695, n_696, n_697, n_698, n_699 : std_logic;
  signal n_700, n_701, n_702, n_703, n_704 : std_logic;
  signal n_705, n_706, n_707, n_708, n_739 : std_logic;
  signal n_742, n_748, n_754, n_760, n_766 : std_logic;
  signal n_772, n_778, n_784, n_790, n_796 : std_logic;
  signal n_802, n_808, n_814, n_820, n_826 : std_logic;
  signal n_832, n_838, n_844, n_850, n_856 : std_logic;
  signal n_862, n_868, n_874, n_880, n_886 : std_logic;
  signal n_892, n_898, n_904, n_910, n_916 : std_logic;
  signal n_922, n_928, n_934, n_940, n_946 : std_logic;
  signal n_952, n_958, n_964, n_970, n_976 : std_logic;
  signal n_982, n_988, n_994, n_1000, n_1006 : std_logic;
  signal n_1012, n_1018, n_1024, n_1030, n_1036 : std_logic;
  signal n_1042, n_1048, n_1054, n_1060, n_1066 : std_logic;
  signal n_1072, n_1078, n_1084, n_1090, n_1096 : std_logic;
  signal n_1102, n_1108, n_1114, n_1120, n_1126 : std_logic;
  signal n_1132, n_1138, n_1144, n_1150, n_1156 : std_logic;
  signal n_1162, n_1168, n_1174, n_1180, n_1186 : std_logic;
  signal n_1192, n_1198, n_1204, n_1210, n_1216 : std_logic;
  signal n_1222, n_1228, n_1234, n_1240, n_1246 : std_logic;
  signal n_1252, n_1258, n_1264, n_1270, n_1276 : std_logic;
  signal n_1282, n_1288, n_1294, n_1300, n_1306 : std_logic;
  signal n_1312, n_1318, n_1324, n_1330, n_1336 : std_logic;
  signal n_1342, n_1348, n_1354, n_1360, n_1366 : std_logic;
  signal n_1372, n_1378, n_1384, n_1390, n_1396 : std_logic;
  signal n_1402, n_1408, n_1414, n_1420, n_1426 : std_logic;
  signal n_1432, n_1438, n_1444, n_1450, n_1456 : std_logic;
  signal n_1462, n_1468, n_1474, n_1480, n_1486 : std_logic;
  signal n_1492, n_1498, n_1504, n_1510, n_1516 : std_logic;
  signal n_1522, n_1528, n_1534, n_1540, n_1546 : std_logic;
  signal n_1552, n_1558, n_1564, n_1570, n_1576 : std_logic;
  signal n_1582, n_1588, n_1594, n_1600, n_1606 : std_logic;
  signal n_1612, n_1618, n_1624, n_1630, n_1636 : std_logic;
  signal n_1642, n_1648, n_1654, n_1660, n_1666 : std_logic;
  signal n_1672, n_1678, n_1684, n_1690, n_1696 : std_logic;
  signal n_1702, n_1708, n_1714, n_1720, n_1726 : std_logic;
  signal n_1732, n_1738, n_1744, n_1750, n_1756 : std_logic;
  signal n_1762, n_1768, n_1774, n_1780, n_1786 : std_logic;
  signal n_1792, n_1798, n_1804, n_1810, n_1816 : std_logic;
  signal n_1820, n_1821 : std_logic;

begin

  framebuffer_buf(116) <= FE_RN_1;
  FE_PHC199_framebuffer_buf_150_3045 : DEL01BWP7T port map(I => FE_PHN171_framebuffer_buf_150_3045, Z => FE_PHN199_framebuffer_buf_150_3045);
  FE_PHC198_framebuffer_buf_101_2996 : DEL01BWP7T port map(I => framebuffer_buf_101_2996, Z => FE_PHN198_framebuffer_buf_101_2996);
  FE_PHC197_framebuffer_buf_106_3001 : DEL01BWP7T port map(I => framebuffer_buf_106_3001, Z => FE_PHN197_framebuffer_buf_106_3001);
  FE_PHC196_framebuffer_buf_79_2974 : DEL01BWP7T port map(I => FE_PHN196_framebuffer_buf_79_2974, Z => framebuffer_buf_79_2974);
  FE_PHC195_framebuffer_buf_126_3021 : DEL01BWP7T port map(I => framebuffer_buf_126_3021, Z => FE_PHN195_framebuffer_buf_126_3021);
  FE_PHC194_framebuffer_buf_118_3013 : DEL01BWP7T port map(I => framebuffer_buf_118_3013, Z => FE_PHN194_framebuffer_buf_118_3013);
  FE_PHC193_framebuffer_buf_80_2975 : DEL01BWP7T port map(I => FE_PHN174_framebuffer_buf_80_2975, Z => FE_PHN193_framebuffer_buf_80_2975);
  FE_PHC192_framebuffer_buf_133_3028 : DEL01BWP7T port map(I => FE_PHN192_framebuffer_buf_133_3028, Z => FE_PHN175_framebuffer_buf_133_3028);
  FE_PHC191_framebuffer_buf_128_3023 : DEL01BWP7T port map(I => FE_PHN191_framebuffer_buf_128_3023, Z => FE_PHN172_framebuffer_buf_128_3023);
  FE_PHC190_framebuffer_buf_154_3049 : DEL01BWP7T port map(I => FE_PHN155_framebuffer_buf_154_3049, Z => FE_PHN190_framebuffer_buf_154_3049);
  FE_PHC189_framebuffer_buf_155_3050 : DEL01BWP7T port map(I => FE_PHN189_framebuffer_buf_155_3050, Z => FE_PHN177_framebuffer_buf_155_3050);
  FE_PHC188_calc_buf_out_2_2873 : DEL01BWP7T port map(I => FE_PHN162_calc_buf_out_2_2873, Z => FE_PHN188_calc_buf_out_2_2873);
  FE_PHC187_framebuffer_buf_93_2988 : DEL01BWP7T port map(I => FE_PHN167_framebuffer_buf_93_2988, Z => FE_PHN187_framebuffer_buf_93_2988);
  FE_PHC186_calc_buf_out_8_2879 : DEL01BWP7T port map(I => FE_PHN176_calc_buf_out_8_2879, Z => FE_PHN186_calc_buf_out_8_2879);
  FE_PHC185_framebuffer_buf_24_2919 : DEL2BWP7T port map(I => framebuffer_buf_24_2919, Z => FE_PHN185_framebuffer_buf_24_2919);
  FE_PHC184_framebuffer_buf_106_3001 : CKBD0BWP7T port map(I => FE_PHN197_framebuffer_buf_106_3001, Z => FE_PHN184_framebuffer_buf_106_3001);
  FE_PHC183_framebuffer_buf_101_2996 : CKBD0BWP7T port map(I => FE_PHN198_framebuffer_buf_101_2996, Z => FE_PHN183_framebuffer_buf_101_2996);
  FE_PHC182_framebuffer_buf_131_3026 : DEL0BWP7T port map(I => framebuffer_buf_131_3026, Z => FE_PHN182_framebuffer_buf_131_3026);
  FE_PHC181_framebuffer_buf_104_2999 : DEL0BWP7T port map(I => framebuffer_buf_104_2999, Z => FE_PHN181_framebuffer_buf_104_2999);
  FE_PHC180_framebuffer_buf_119_3014 : DEL0BWP7T port map(I => FE_PHN180_framebuffer_buf_119_3014, Z => framebuffer_buf_119_3014);
  FE_PHC179_framebuffer_buf_89_2984 : DEL1BWP7T port map(I => framebuffer_buf_89_2984, Z => FE_PHN179_framebuffer_buf_89_2984);
  FE_PHC178_framebuffer_buf_4_2899 : DEL0BWP7T port map(I => framebuffer_buf_4_2899, Z => FE_PHN178_framebuffer_buf_4_2899);
  FE_PHC177_framebuffer_buf_155_3050 : CKBD0BWP7T port map(I => FE_PHN177_framebuffer_buf_155_3050, Z => framebuffer_buf_155_3050);
  FE_PHC176_calc_buf_out_8_2879 : CKBD0BWP7T port map(I => calc_buf_out_8_2879, Z => FE_PHN176_calc_buf_out_8_2879);
  FE_PHC175_framebuffer_buf_133_3028 : CKBD0BWP7T port map(I => FE_PHN175_framebuffer_buf_133_3028, Z => framebuffer_buf_133_3028);
  FE_PHC174_framebuffer_buf_80_2975 : CKBD0BWP7T port map(I => framebuffer_buf_80_2975, Z => FE_PHN174_framebuffer_buf_80_2975);
  FE_PHC173_framebuffer_buf_127_3022 : DEL1BWP7T port map(I => framebuffer_buf_127_3022, Z => FE_PHN173_framebuffer_buf_127_3022);
  FE_PHC172_framebuffer_buf_128_3023 : CKBD0BWP7T port map(I => FE_PHN172_framebuffer_buf_128_3023, Z => framebuffer_buf_128_3023);
  FE_PHC171_framebuffer_buf_150_3045 : CKBD0BWP7T port map(I => framebuffer_buf_150_3045, Z => FE_PHN171_framebuffer_buf_150_3045);
  FE_PHC170_framebuffer_buf_126_3021 : CKBD0BWP7T port map(I => FE_PHN195_framebuffer_buf_126_3021, Z => FE_PHN170_framebuffer_buf_126_3021);
  FE_PHC169_framebuffer_buf_71_2966 : DEL0BWP7T port map(I => FE_PHN169_framebuffer_buf_71_2966, Z => framebuffer_buf_71_2966);
  FE_PHC168_framebuffer_buf_146_3041 : DEL0BWP7T port map(I => framebuffer_buf_146_3041, Z => FE_PHN168_framebuffer_buf_146_3041);
  FE_PHC167_framebuffer_buf_93_2988 : CKBD0BWP7T port map(I => framebuffer_buf_93_2988, Z => FE_PHN167_framebuffer_buf_93_2988);
  FE_PHC166_framebuffer_buf_5_2900 : DEL0BWP7T port map(I => framebuffer_buf_5_2900, Z => FE_PHN166_framebuffer_buf_5_2900);
  FE_PHC165_framebuffer_buf_152_3047 : DEL0BWP7T port map(I => framebuffer_buf_152_3047, Z => FE_PHN165_framebuffer_buf_152_3047);
  FE_PHC164_calc_buf_out_13_2884 : DEL1BWP7T port map(I => calc_buf_out_13_2884, Z => FE_PHN164_calc_buf_out_13_2884);
  FE_PHC163_framebuffer_buf_84_2979 : DEL0BWP7T port map(I => framebuffer_buf_84_2979, Z => FE_PHN163_framebuffer_buf_84_2979);
  FE_PHC162_calc_buf_out_2_2873 : CKBD0BWP7T port map(I => calc_buf_out_2_2873, Z => FE_PHN162_calc_buf_out_2_2873);
  FE_PHC161_framebuffer_buf_99_2994 : DEL0BWP7T port map(I => framebuffer_buf_99_2994, Z => FE_PHN161_framebuffer_buf_99_2994);
  FE_PHC160_framebuffer_buf_40_2935 : DEL0BWP7T port map(I => framebuffer_buf_40_2935, Z => FE_PHN160_framebuffer_buf_40_2935);
  FE_PHC159_framebuffer_buf_122_3017 : DEL1BWP7T port map(I => framebuffer_buf_122_3017, Z => FE_PHN159_framebuffer_buf_122_3017);
  FE_PHC158_framebuffer_buf_86_2981 : CKBD3BWP7T port map(I => framebuffer_buf_86_2981, Z => FE_PHN158_framebuffer_buf_86_2981);
  FE_PHC157_framebuffer_buf_79_2974 : CKBD0BWP7T port map(I => framebuffer_buf_79_2974, Z => FE_PHN157_framebuffer_buf_79_2974);
  FE_PHC156_framebuffer_buf_103_2998 : DEL0BWP7T port map(I => framebuffer_buf_103_2998, Z => FE_PHN156_framebuffer_buf_103_2998);
  FE_PHC155_framebuffer_buf_154_3049 : CKBD0BWP7T port map(I => framebuffer_buf_154_3049, Z => FE_PHN155_framebuffer_buf_154_3049);
  FE_PHC154_framebuffer_buf_70_2965 : DEL0BWP7T port map(I => framebuffer_buf_70_2965, Z => FE_PHN154_framebuffer_buf_70_2965);
  FE_PHC153_framebuffer_buf_53_2948 : DEL0BWP7T port map(I => framebuffer_buf_53_2948, Z => FE_PHN153_framebuffer_buf_53_2948);
  FE_PHC152_calc_buf_out_21_2892 : DEL0BWP7T port map(I => calc_buf_out_21_2892, Z => FE_PHN152_calc_buf_out_21_2892);
  FE_PHC151_framebuffer_buf_120_3015 : DEL0BWP7T port map(I => FE_PHN151_framebuffer_buf_120_3015, Z => framebuffer_buf_120_3015);
  FE_PHC150_framebuffer_buf_118_3013 : CKBD0BWP7T port map(I => FE_PHN194_framebuffer_buf_118_3013, Z => FE_PHN150_framebuffer_buf_118_3013);
  FE_PHC149_framebuffer_buf_49_2944 : DEL0BWP7T port map(I => framebuffer_buf_49_2944, Z => FE_PHN149_framebuffer_buf_49_2944);
  FE_PHC148_framebuffer_buf_157_3052 : DEL0BWP7T port map(I => FE_PHN148_framebuffer_buf_157_3052, Z => framebuffer_buf_157_3052);
  FE_PHC147_framebuffer_buf_156_3051 : DEL0BWP7T port map(I => framebuffer_buf_156_3051, Z => FE_PHN147_framebuffer_buf_156_3051);
  FE_PHC146_framebuffer_buf_55_2950 : DEL1BWP7T port map(I => FE_PHN146_framebuffer_buf_55_2950, Z => framebuffer_buf_55_2950);
  FE_PHC145_framebuffer_buf_47_2942 : DEL1BWP7T port map(I => framebuffer_buf_47_2942, Z => FE_PHN145_framebuffer_buf_47_2942);
  FE_PHC144_framebuffer_buf_44_2939 : DEL1BWP7T port map(I => framebuffer_buf_44_2939, Z => FE_PHN144_framebuffer_buf_44_2939);
  FE_PHC143_framebuffer_buf_37_2932 : DEL1BWP7T port map(I => FE_PHN143_framebuffer_buf_37_2932, Z => framebuffer_buf_37_2932);
  FE_PHC142_framebuffer_buf_78_2973 : DEL0BWP7T port map(I => framebuffer_buf_78_2973, Z => FE_PHN142_framebuffer_buf_78_2973);
  FE_PHC141_framebuffer_buf_132_3027 : DEL0BWP7T port map(I => FE_PHN141_framebuffer_buf_132_3027, Z => framebuffer_buf_132_3027);
  FE_PHC140_framebuffer_buf_43_2938 : DEL0BWP7T port map(I => framebuffer_buf_43_2938, Z => FE_PHN140_framebuffer_buf_43_2938);
  FE_PHC139_framebuffer_buf_143_3038 : DEL0BWP7T port map(I => framebuffer_buf_143_3038, Z => FE_PHN139_framebuffer_buf_143_3038);
  FE_PHC138_framebuffer_buf_88_2983 : DEL01BWP7T port map(I => framebuffer_buf_88_2983, Z => FE_PHN138_framebuffer_buf_88_2983);
  FE_PHC137_framebuffer_buf_129_3024 : DEL0BWP7T port map(I => FE_PHN137_framebuffer_buf_129_3024, Z => framebuffer_buf_129_3024);
  FE_PHC136_framebuffer_buf_12_2907 : DEL0BWP7T port map(I => framebuffer_buf_12_2907, Z => FE_PHN136_framebuffer_buf_12_2907);
  FE_PHC135_calc_buf_out_18_2889 : DEL0BWP7T port map(I => calc_buf_out_18_2889, Z => FE_PHN135_calc_buf_out_18_2889);
  FE_PHC134_framebuffer_buf_13_2908 : DEL0BWP7T port map(I => framebuffer_buf_13_2908, Z => FE_PHN134_framebuffer_buf_13_2908);
  FE_PHC133_framebuffer_buf_14_2909 : DEL0BWP7T port map(I => framebuffer_buf_14_2909, Z => FE_PHN133_framebuffer_buf_14_2909);
  FE_PHC132_framebuffer_buf_124_3019 : DEL0BWP7T port map(I => framebuffer_buf_124_3019, Z => FE_PHN132_framebuffer_buf_124_3019);
  FE_PHC131_framebuffer_buf_72_2967 : DEL0BWP7T port map(I => framebuffer_buf_72_2967, Z => FE_PHN131_framebuffer_buf_72_2967);
  FE_PHC130_framebuffer_buf_83_2978 : DEL0BWP7T port map(I => framebuffer_buf_83_2978, Z => FE_PHN130_framebuffer_buf_83_2978);
  FE_PHC129_framebuffer_buf_96_2991 : DEL0BWP7T port map(I => framebuffer_buf_96_2991, Z => FE_PHN129_framebuffer_buf_96_2991);
  FE_PHC128_framebuffer_buf_62_2957 : DEL0BWP7T port map(I => framebuffer_buf_62_2957, Z => FE_PHN128_framebuffer_buf_62_2957);
  FE_PHC127_framebuffer_buf_142_3037 : DEL0BWP7T port map(I => framebuffer_buf_142_3037, Z => FE_PHN127_framebuffer_buf_142_3037);
  FE_PHC126_framebuffer_buf_153_3048 : DEL0BWP7T port map(I => framebuffer_buf_153_3048, Z => FE_PHN126_framebuffer_buf_153_3048);
  FE_PHC125_framebuffer_buf_149_3044 : DEL0BWP7T port map(I => FE_PHN125_framebuffer_buf_149_3044, Z => framebuffer_buf_149_3044);
  FE_PHC124_framebuffer_buf_76_2971 : DEL0BWP7T port map(I => framebuffer_buf_76_2971, Z => FE_PHN124_framebuffer_buf_76_2971);
  FE_PHC123_framebuffer_buf_111_3006 : DEL0BWP7T port map(I => framebuffer_buf_111_3006, Z => FE_PHN123_framebuffer_buf_111_3006);
  FE_PHC122_framebuffer_buf_112_3007 : DEL0BWP7T port map(I => framebuffer_buf_112_3007, Z => FE_PHN122_framebuffer_buf_112_3007);
  FE_PHC121_framebuffer_buf_134_3029 : DEL0BWP7T port map(I => framebuffer_buf_134_3029, Z => FE_PHN121_framebuffer_buf_134_3029);
  FE_PHC120_framebuffer_buf_147_3042 : DEL0BWP7T port map(I => framebuffer_buf_147_3042, Z => FE_PHN120_framebuffer_buf_147_3042);
  FE_PHC119_framebuffer_buf_130_3025 : DEL0BWP7T port map(I => FE_PHN119_framebuffer_buf_130_3025, Z => framebuffer_buf_130_3025);
  FE_PHC118_framebuffer_buf_114_3009 : DEL0BWP7T port map(I => framebuffer_buf_114_3009, Z => FE_PHN118_framebuffer_buf_114_3009);
  FE_PHC117_framebuffer_buf_27_2922 : DEL0BWP7T port map(I => framebuffer_buf_27_2922, Z => FE_PHN117_framebuffer_buf_27_2922);
  FE_PHC116_framebuffer_buf_144_3039 : BUFFD3BWP7T port map(I => framebuffer_buf_144_3039, Z => FE_PHN116_framebuffer_buf_144_3039);
  FE_PHC115_framebuffer_buf_105_3000 : DEL0BWP7T port map(I => framebuffer_buf_105_3000, Z => FE_PHN115_framebuffer_buf_105_3000);
  FE_PHC114_framebuffer_buf_113_3008 : DEL0BWP7T port map(I => FE_PHN114_framebuffer_buf_113_3008, Z => framebuffer_buf_113_3008);
  FE_PHC113_framebuffer_buf_98_2993 : DEL0BWP7T port map(I => framebuffer_buf_98_2993, Z => FE_PHN113_framebuffer_buf_98_2993);
  FE_PHC112_framebuffer_buf_33_2928 : DEL0BWP7T port map(I => framebuffer_buf_33_2928, Z => FE_PHN112_framebuffer_buf_33_2928);
  FE_PHC111_framebuffer_buf_6_2901 : DEL0BWP7T port map(I => framebuffer_buf_6_2901, Z => FE_PHN111_framebuffer_buf_6_2901);
  FE_PHC110_framebuffer_buf_87_2982 : DEL0BWP7T port map(I => framebuffer_buf_87_2982, Z => FE_PHN110_framebuffer_buf_87_2982);
  FE_PHC109_framebuffer_buf_17_2912 : DEL0BWP7T port map(I => FE_PHN109_framebuffer_buf_17_2912, Z => framebuffer_buf_17_2912);
  FE_PHC108_framebuffer_buf_63_2958 : DEL0BWP7T port map(I => framebuffer_buf_63_2958, Z => FE_PHN108_framebuffer_buf_63_2958);
  FE_PHC107_framebuffer_buf_67_2962 : BUFFD3BWP7T port map(I => framebuffer_buf_67_2962, Z => FE_PHN107_framebuffer_buf_67_2962);
  FE_PHC106_framebuffer_buf_46_2941 : DEL0BWP7T port map(I => framebuffer_buf_46_2941, Z => FE_PHN106_framebuffer_buf_46_2941);
  FE_PHC105_framebuffer_buf_77_2972 : DEL0BWP7T port map(I => framebuffer_buf_77_2972, Z => FE_PHN105_framebuffer_buf_77_2972);
  FE_PHC104_framebuffer_buf_65_2960 : DEL0BWP7T port map(I => framebuffer_buf_65_2960, Z => FE_PHN104_framebuffer_buf_65_2960);
  FE_PHC103_framebuffer_buf_110_3005 : DEL0BWP7T port map(I => framebuffer_buf_110_3005, Z => FE_PHN103_framebuffer_buf_110_3005);
  FE_PHC102_framebuffer_buf_141_3036 : DEL0BWP7T port map(I => framebuffer_buf_141_3036, Z => FE_PHN102_framebuffer_buf_141_3036);
  FE_PHC101_framebuffer_buf_8_2903 : DEL0BWP7T port map(I => framebuffer_buf_8_2903, Z => FE_PHN101_framebuffer_buf_8_2903);
  FE_PHC100_framebuffer_buf_42_2937 : DEL0BWP7T port map(I => framebuffer_buf_42_2937, Z => FE_PHN100_framebuffer_buf_42_2937);
  FE_PHC99_framebuffer_buf_52_2947 : DEL0BWP7T port map(I => framebuffer_buf_52_2947, Z => FE_PHN99_framebuffer_buf_52_2947);
  FE_PHC98_framebuffer_buf_15_2910 : DEL0BWP7T port map(I => framebuffer_buf_15_2910, Z => FE_PHN98_framebuffer_buf_15_2910);
  FE_PHC97_framebuffer_buf_137_3032 : DEL0BWP7T port map(I => framebuffer_buf_137_3032, Z => FE_PHN97_framebuffer_buf_137_3032);
  FE_PHC96_framebuffer_buf_39_2934 : DEL0BWP7T port map(I => framebuffer_buf_39_2934, Z => FE_PHN96_framebuffer_buf_39_2934);
  FE_PHC95_framebuffer_buf_19_2914 : DEL0BWP7T port map(I => framebuffer_buf_19_2914, Z => FE_PHN95_framebuffer_buf_19_2914);
  FE_PHC94_calc_buf_out_19_2890 : DEL0BWP7T port map(I => calc_buf_out_19_2890, Z => FE_PHN94_calc_buf_out_19_2890);
  FE_PHC93_framebuffer_buf_75_2970 : DEL0BWP7T port map(I => framebuffer_buf_75_2970, Z => FE_PHN93_framebuffer_buf_75_2970);
  FE_PHC92_framebuffer_buf_145_3040 : DEL0BWP7T port map(I => framebuffer_buf_145_3040, Z => FE_PHN92_framebuffer_buf_145_3040);
  FE_PHC91_framebuffer_buf_51_2946 : DEL0BWP7T port map(I => framebuffer_buf_51_2946, Z => FE_PHN91_framebuffer_buf_51_2946);
  FE_PHC90_framebuffer_buf_34_2929 : DEL0BWP7T port map(I => framebuffer_buf_34_2929, Z => FE_PHN90_framebuffer_buf_34_2929);
  FE_PHC89_framebuffer_buf_69_2964 : DEL0BWP7T port map(I => framebuffer_buf_69_2964, Z => FE_PHN89_framebuffer_buf_69_2964);
  FE_PHC88_framebuffer_buf_48_2943 : DEL0BWP7T port map(I => framebuffer_buf_48_2943, Z => FE_PHN88_framebuffer_buf_48_2943);
  FE_PHC87_framebuffer_buf_58_2953 : DEL0BWP7T port map(I => FE_PHN87_framebuffer_buf_58_2953, Z => framebuffer_buf_58_2953);
  FE_PHC86_framebuffer_buf_25_2920 : DEL0BWP7T port map(I => framebuffer_buf_25_2920, Z => FE_PHN86_framebuffer_buf_25_2920);
  FE_PHC85_framebuffer_buf_16_2911 : DEL0BWP7T port map(I => framebuffer_buf_16_2911, Z => FE_PHN85_framebuffer_buf_16_2911);
  FE_PHC84_calc_buf_out_7_2878 : DEL0BWP7T port map(I => calc_buf_out_7_2878, Z => FE_PHN84_calc_buf_out_7_2878);
  FE_PHC83_calc_buf_out_6_2877 : DEL0BWP7T port map(I => calc_buf_out_6_2877, Z => FE_PHN83_calc_buf_out_6_2877);
  FE_PHC82_framebuffer_buf_18_2913 : DEL0BWP7T port map(I => framebuffer_buf_18_2913, Z => FE_PHN82_framebuffer_buf_18_2913);
  FE_PHC81_framebuffer_buf_140_3035 : DEL0BWP7T port map(I => framebuffer_buf_140_3035, Z => FE_PHN81_framebuffer_buf_140_3035);
  FE_PHC80_framebuffer_buf_64_2959 : DEL0BWP7T port map(I => framebuffer_buf_64_2959, Z => FE_PHN80_framebuffer_buf_64_2959);
  FE_PHC79_framebuffer_buf_95_2990 : DEL0BWP7T port map(I => framebuffer_buf_95_2990, Z => FE_PHN79_framebuffer_buf_95_2990);
  FE_PHC78_framebuffer_buf_109_3004 : DEL0BWP7T port map(I => framebuffer_buf_109_3004, Z => FE_PHN78_framebuffer_buf_109_3004);
  FE_PHC77_framebuffer_buf_148_3043 : DEL0BWP7T port map(I => framebuffer_buf_148_3043, Z => FE_PHN77_framebuffer_buf_148_3043);
  FE_PHC76_framebuffer_buf_22_2917 : DEL0BWP7T port map(I => framebuffer_buf_22_2917, Z => FE_PHN76_framebuffer_buf_22_2917);
  FE_PHC75_calc_buf_out_14_2885 : DEL0BWP7T port map(I => calc_buf_out_14_2885, Z => FE_PHN75_calc_buf_out_14_2885);
  FE_PHC74_framebuffer_buf_68_2963 : DEL0BWP7T port map(I => framebuffer_buf_68_2963, Z => FE_PHN74_framebuffer_buf_68_2963);
  FE_PHC73_framebuffer_buf_151_3046 : DEL0BWP7T port map(I => framebuffer_buf_151_3046, Z => FE_PHN73_framebuffer_buf_151_3046);
  FE_PHC72_framebuffer_buf_60_2955 : DEL0BWP7T port map(I => framebuffer_buf_60_2955, Z => FE_PHN72_framebuffer_buf_60_2955);
  FE_PHC71_framebuffer_buf_136_3031 : DEL0BWP7T port map(I => FE_PHN71_framebuffer_buf_136_3031, Z => framebuffer_buf_136_3031);
  FE_PHC70_framebuffer_buf_36_2931 : DEL0BWP7T port map(I => framebuffer_buf_36_2931, Z => FE_PHN70_framebuffer_buf_36_2931);
  FE_PHC69_framebuffer_buf_28_2923 : DEL0BWP7T port map(I => FE_PHN69_framebuffer_buf_28_2923, Z => framebuffer_buf_28_2923);
  FE_PHC68_calc_buf_out_10_2881 : DEL0BWP7T port map(I => FE_PHN68_calc_buf_out_10_2881, Z => calc_buf_out_10_2881);
  FE_PHC67_framebuffer_buf_21_2916 : DEL0BWP7T port map(I => framebuffer_buf_21_2916, Z => FE_PHN67_framebuffer_buf_21_2916);
  FE_PHC66_framebuffer_buf_41_2936 : DEL0BWP7T port map(I => FE_PHN66_framebuffer_buf_41_2936, Z => framebuffer_buf_41_2936);
  FE_PHC65_framebuffer_buf_56_2951 : DEL0BWP7T port map(I => framebuffer_buf_56_2951, Z => FE_PHN65_framebuffer_buf_56_2951);
  FE_PHC64_calc_buf_out_15_2886 : DEL0BWP7T port map(I => calc_buf_out_15_2886, Z => FE_PHN64_calc_buf_out_15_2886);
  FE_PHC63_framebuffer_buf_73_2968 : DEL0BWP7T port map(I => framebuffer_buf_73_2968, Z => FE_PHN63_framebuffer_buf_73_2968);
  FE_PHC62_framebuffer_buf_123_3018 : DEL0BWP7T port map(I => FE_PHN62_framebuffer_buf_123_3018, Z => framebuffer_buf_123_3018);
  FE_PHC61_framebuffer_buf_108_3003 : DEL0BWP7T port map(I => framebuffer_buf_108_3003, Z => FE_PHN61_framebuffer_buf_108_3003);
  FE_PHC60_framebuffer_buf_102_2997 : DEL0BWP7T port map(I => framebuffer_buf_102_2997, Z => FE_PHN60_framebuffer_buf_102_2997);
  FE_PHC59_framebuffer_buf_139_3034 : DEL0BWP7T port map(I => framebuffer_buf_139_3034, Z => FE_PHN59_framebuffer_buf_139_3034);
  FE_PHC58_framebuffer_buf_94_2989 : DEL0BWP7T port map(I => framebuffer_buf_94_2989, Z => FE_PHN58_framebuffer_buf_94_2989);
  FE_PHC57_framebuffer_buf_35_2930 : DEL0BWP7T port map(I => framebuffer_buf_35_2930, Z => FE_PHN57_framebuffer_buf_35_2930);
  FE_PHC56_framebuffer_buf_138_3033 : DEL0BWP7T port map(I => framebuffer_buf_138_3033, Z => FE_PHN56_framebuffer_buf_138_3033);
  FE_PHC55_framebuffer_buf_97_2992 : DEL0BWP7T port map(I => framebuffer_buf_97_2992, Z => FE_PHN55_framebuffer_buf_97_2992);
  FE_PHC54_framebuffer_buf_115_3010 : DEL0BWP7T port map(I => FE_PHN54_framebuffer_buf_115_3010, Z => framebuffer_buf_115_3010);
  FE_PHC53_framebuffer_buf_11_2906 : DEL0BWP7T port map(I => framebuffer_buf_11_2906, Z => FE_PHN53_framebuffer_buf_11_2906);
  FE_PHC52_framebuffer_buf_45_2940 : DEL0BWP7T port map(I => framebuffer_buf_45_2940, Z => FE_PHN52_framebuffer_buf_45_2940);
  FE_PHC51_framebuffer_buf_50_2945 : DEL0BWP7T port map(I => framebuffer_buf_50_2945, Z => FE_PHN51_framebuffer_buf_50_2945);
  FE_PHC50_framebuffer_buf_135_3030 : DEL0BWP7T port map(I => FE_PHN50_framebuffer_buf_135_3030, Z => framebuffer_buf_135_3030);
  FE_PHC49_calc_buf_out_11_2882 : DEL0BWP7T port map(I => calc_buf_out_11_2882, Z => FE_PHN49_calc_buf_out_11_2882);
  FE_PHC48_framebuffer_buf_66_2961 : DEL0BWP7T port map(I => framebuffer_buf_66_2961, Z => FE_PHN48_framebuffer_buf_66_2961);
  FE_PHC47_framebuffer_buf_74_2969 : DEL0BWP7T port map(I => framebuffer_buf_74_2969, Z => FE_PHN47_framebuffer_buf_74_2969);
  FE_PHC46_framebuffer_buf_125_3020 : DEL0BWP7T port map(I => framebuffer_buf_125_3020, Z => FE_PHN46_framebuffer_buf_125_3020);
  FE_PHC45_framebuffer_buf_9_2904 : DEL0BWP7T port map(I => framebuffer_buf_9_2904, Z => FE_PHN45_framebuffer_buf_9_2904);
  FE_PHC44_framebuffer_buf_31_2926 : DEL0BWP7T port map(I => framebuffer_buf_31_2926, Z => FE_PHN44_framebuffer_buf_31_2926);
  FE_PHC43_framebuffer_buf_1_2896 : DEL0BWP7T port map(I => framebuffer_buf_1_2896, Z => FE_PHN43_framebuffer_buf_1_2896);
  FE_PHC42_framebuffer_buf_107_3002 : DEL0BWP7T port map(I => framebuffer_buf_107_3002, Z => FE_PHN42_framebuffer_buf_107_3002);
  FE_PHC41_framebuffer_buf_26_2921 : DEL0BWP7T port map(I => framebuffer_buf_26_2921, Z => FE_PHN41_framebuffer_buf_26_2921);
  FE_PHC40_framebuffer_buf_0_2895 : DEL0BWP7T port map(I => framebuffer_buf_0_2895, Z => FE_PHN40_framebuffer_buf_0_2895);
  FE_PHC39_framebuffer_buf_54_2949 : DEL0BWP7T port map(I => framebuffer_buf_54_2949, Z => FE_PHN39_framebuffer_buf_54_2949);
  FE_PHC38_framebuffer_buf_10_2905 : DEL0BWP7T port map(I => framebuffer_buf_10_2905, Z => FE_PHN38_framebuffer_buf_10_2905);
  FE_PHC37_calc_buf_out_5_2876 : DEL0BWP7T port map(I => calc_buf_out_5_2876, Z => FE_PHN37_calc_buf_out_5_2876);
  FE_PHC36_framebuffer_buf_23_2918 : DEL0BWP7T port map(I => FE_PHN36_framebuffer_buf_23_2918, Z => framebuffer_buf_23_2918);
  FE_PHC35_framebuffer_buf_38_2933 : DEL0BWP7T port map(I => framebuffer_buf_38_2933, Z => FE_PHN35_framebuffer_buf_38_2933);
  FE_PHC34_framebuffer_buf_32_2927 : DEL0BWP7T port map(I => framebuffer_buf_32_2927, Z => FE_PHN34_framebuffer_buf_32_2927);
  FE_PHC33_framebuffer_buf_121_3016 : DEL0BWP7T port map(I => framebuffer_buf_121_3016, Z => FE_PHN33_framebuffer_buf_121_3016);
  FE_PHC32_calc_buf_out_12_2883 : DEL0BWP7T port map(I => calc_buf_out_12_2883, Z => FE_PHN32_calc_buf_out_12_2883);
  FE_PHC31_calc_buf_out_22_2893 : DEL0BWP7T port map(I => calc_buf_out_22_2893, Z => FE_PHN31_calc_buf_out_22_2893);
  FE_PHC30_calc_buf_out_4_2875 : DEL0BWP7T port map(I => calc_buf_out_4_2875, Z => FE_PHN30_calc_buf_out_4_2875);
  FE_PHC29_framebuffer_buf_92_2987 : DEL0BWP7T port map(I => framebuffer_buf_92_2987, Z => FE_PHN29_framebuffer_buf_92_2987);
  FE_PHC28_calc_buf_out_3_2874 : DEL0BWP7T port map(I => calc_buf_out_3_2874, Z => FE_PHN28_calc_buf_out_3_2874);
  FE_PHC27_framebuffer_buf_57_2952 : DEL0BWP7T port map(I => framebuffer_buf_57_2952, Z => FE_PHN27_framebuffer_buf_57_2952);
  FE_PHC26_framebuffer_buf_100_2995 : DEL0BWP7T port map(I => framebuffer_buf_100_2995, Z => FE_PHN26_framebuffer_buf_100_2995);
  FE_PHC25_calc_buf_out_20_2891 : DEL0BWP7T port map(I => calc_buf_out_20_2891, Z => FE_PHN25_calc_buf_out_20_2891);
  FE_PHC24_framebuffer_buf_61_2956 : DEL0BWP7T port map(I => framebuffer_buf_61_2956, Z => FE_PHN24_framebuffer_buf_61_2956);
  FE_PHC23_calc_buf_out_23_2894 : DEL0BWP7T port map(I => calc_buf_out_23_2894, Z => FE_PHN23_calc_buf_out_23_2894);
  FE_PHC22_framebuffer_buf_30_2925 : DEL0BWP7T port map(I => framebuffer_buf_30_2925, Z => FE_PHN22_framebuffer_buf_30_2925);
  FE_PHC21_framebuffer_buf_2_2897 : DEL0BWP7T port map(I => framebuffer_buf_2_2897, Z => FE_PHN21_framebuffer_buf_2_2897);
  FE_PHC20_framebuffer_buf_29_2924 : DEL0BWP7T port map(I => framebuffer_buf_29_2924, Z => FE_PHN20_framebuffer_buf_29_2924);
  FE_PHC19_framebuffer_buf_3_2898 : DEL0BWP7T port map(I => FE_PHN19_framebuffer_buf_3_2898, Z => framebuffer_buf_3_2898);
  FE_PHC18_framebuffer_buf_20_2915 : DEL0BWP7T port map(I => framebuffer_buf_20_2915, Z => FE_PHN18_framebuffer_buf_20_2915);
  FE_PHC17_calc_buf_out_17_2888 : DEL0BWP7T port map(I => calc_buf_out_17_2888, Z => FE_PHN17_calc_buf_out_17_2888);
  FE_PHC16_calc_buf_out_9_2880 : DEL0BWP7T port map(I => FE_PHN16_calc_buf_out_9_2880, Z => calc_buf_out_9_2880);
  FE_PHC15_calc_buf_out_16_2887 : DEL0BWP7T port map(I => calc_buf_out_16_2887, Z => FE_PHN15_calc_buf_out_16_2887);
  FE_PHC14_calc_buf_out_1_2872 : DEL0BWP7T port map(I => calc_buf_out_1_2872, Z => FE_PHN14_calc_buf_out_1_2872);
  FE_PHC13_calc_buf_out_0_2871 : DEL0BWP7T port map(I => calc_buf_out_0_2871, Z => FE_PHN13_calc_buf_out_0_2871);
  FE_PHC12_framebuffer_buf_90_2985 : DEL01BWP7T port map(I => framebuffer_buf_90_2985, Z => FE_PHN12_framebuffer_buf_90_2985);
  FE_PHC11_framebuffer_buf_91_2986 : DEL01BWP7T port map(I => framebuffer_buf_91_2986, Z => FE_PHN11_framebuffer_buf_91_2986);
  FE_PHC10_framebuffer_buf_82_2977 : DEL01BWP7T port map(I => framebuffer_buf_82_2977, Z => FE_PHN10_framebuffer_buf_82_2977);
  FE_PHC9_framebuffer_buf_7_2902 : CKBD0BWP7T port map(I => framebuffer_buf_7_2902, Z => FE_PHN9_framebuffer_buf_7_2902);
  FE_PHC8_framebuffer_buf_85_2980 : CKBD0BWP7T port map(I => FE_PHN8_framebuffer_buf_85_2980, Z => framebuffer_buf_85_2980);
  FE_PHC7_framebuffer_buf_81_2976 : CKBD0BWP7T port map(I => framebuffer_buf_81_2976, Z => FE_PHN7_framebuffer_buf_81_2976);
  FE_PHC6_framebuffer_buf_59_2954 : CKBD0BWP7T port map(I => framebuffer_buf_59_2954, Z => FE_PHN6_framebuffer_buf_59_2954);
  FE_OFC5_framebuffer_buf_116 : BUFFD5BWP7T port map(I => framebuffer_buf(116), Z => framebuffer_buf(117));
  FE_OFC4_framebuffer_buf_116 : BUFFD5BWP7T port map(I => FE_OFN4_framebuffer_buf_116, Z => FE_RN_1);
  FE_OFC3_n_0 : BUFFD2BWP7T port map(I => FE_OFN1_n_0, Z => FE_OFN3_n_0);
  FE_OFC2_n_0 : INVD1BWP7T port map(I => FE_OFN0_n_0, ZN => FE_OFN2_n_0);
  FE_OFC1_n_0 : CKND2BWP7T port map(I => FE_OFN0_n_0, ZN => FE_OFN1_n_0);
  FE_OFC0_n_0 : INVD1BWP7T port map(I => n_0, ZN => FE_OFN0_n_0);
  CTS_ccl_a_BUF_clk_G0_L2_3 : CKBD12BWP7T port map(I => CTS_16, Z => CTS_15);
  CTS_ccl_a_BUF_clk_G0_L2_2 : CKBD12BWP7T port map(I => CTS_16, Z => CTS_14);
  CTS_ccl_a_BUF_clk_G0_L2_1 : CKBD12BWP7T port map(I => CTS_16, Z => CTS_13);
  CTS_ccl_a_BUF_clk_G0_L1_1 : CKBD8BWP7T port map(I => clk, Z => CTS_16);
  new_sqi_address_reg_12 : LHQD1BWP7T port map(D => n_682, E => n_681, Q => new_sqi_address(12));
  g24617 : ND2D0BWP7T port map(A1 => n_680, A2 => n_372, ZN => n_682);
  new_sqi_address_reg_13 : LHQD1BWP7T port map(D => n_679, E => n_681, Q => new_sqi_address(13));
  new_sqi_address_reg_11 : LHQD1BWP7T port map(D => n_678, E => n_681, Q => new_sqi_address(11));
  g24628 : AOI211D0BWP7T port map(A1 => n_272, A2 => n_258, B => n_676, C => n_367, ZN => n_680);
  new_sqi_address_reg_14 : LHQD1BWP7T port map(D => n_675, E => n_681, Q => new_sqi_address(14));
  g24613 : ND3D0BWP7T port map(A1 => n_677, A2 => n_667, A3 => n_674, ZN => n_679);
  g24625 : ND4D0BWP7T port map(A1 => n_670, A2 => n_422, A3 => n_159, A4 => n_210, ZN => n_678);
  g24618 : AOI31D0BWP7T port map(A1 => n_668, A2 => n_363, A3 => n_6, B => n_671, ZN => n_677);
  g24686 : OAI31D0BWP7T port map(A1 => counter(6), A2 => n_369, A3 => n_377, B => n_672, ZN => n_676);
  g24627 : ND4D0BWP7T port map(A1 => n_669, A2 => n_674, A3 => n_408, A4 => n_368, ZN => n_675);
  new_sqi_address_reg_10 : LHQD1BWP7T port map(D => n_666, E => n_681, Q => new_sqi_address(10));
  g24785 : NR4D0BWP7T port map(A1 => n_543, A2 => n_420, A3 => n_365, A4 => n_182, ZN => n_672);
  g24626 : IND4D0BWP7T port map(A1 => n_572, B1 => n_190, B2 => n_184, B3 => n_202, ZN => n_671);
  g24832 : AOI31D0BWP7T port map(A1 => n_209, A2 => n_418, A3 => n_183, B => n_664, ZN => n_670);
  new_sqi_address_reg_9 : LHQD1BWP7T port map(D => n_665, E => n_681, Q => new_sqi_address(9));
  g24830 : AOI211D0BWP7T port map(A1 => n_668, A2 => n_59, B => n_505, C => n_198, ZN => n_669);
  g24999 : AOI222D0BWP7T port map(A1 => n_484, A2 => counter(7), B1 => n_373, B2 => n_504, C1 => n_370, C2 => counter(7), ZN => n_667);
  g24784 : ND4D0BWP7T port map(A1 => n_503, A2 => n_179, A3 => n_270, A4 => n_188, ZN => n_666);
  g25046 : OAI211D0BWP7T port map(A1 => n_327, A2 => n_232, B => n_489, C => n_117, ZN => n_665);
  g24979 : MOAI22D0BWP7T port map(A1 => n_485, A2 => counter(5), B1 => n_488, B2 => sqi_address(11), ZN => n_664);
  g24926 : MOAI22D0BWP7T port map(A1 => n_597, A2 => n_625, B1 => n_595, B2 => FE_PHN121_framebuffer_buf_134_3029, ZN => n_662);
  g24887 : MOAI22D0BWP7T port map(A1 => n_659, A2 => n_653, B1 => n_658, B2 => FE_PHN97_framebuffer_buf_137_3032, ZN => n_661);
  g24888 : MOAI22D0BWP7T port map(A1 => n_659, A2 => n_650, B1 => n_658, B2 => FE_PHN56_framebuffer_buf_138_3033, ZN => n_660);
  g24889 : MOAI22D0BWP7T port map(A1 => n_659, A2 => n_648, B1 => n_658, B2 => FE_PHN59_framebuffer_buf_139_3034, ZN => n_657);
  g24890 : MOAI22D0BWP7T port map(A1 => n_654, A2 => n_641, B1 => n_652, B2 => FE_PHN128_framebuffer_buf_62_2957, ZN => n_656);
  g24891 : MOAI22D0BWP7T port map(A1 => n_654, A2 => n_653, B1 => n_652, B2 => FE_PHN108_framebuffer_buf_63_2958, ZN => n_655);
  g24892 : MOAI22D0BWP7T port map(A1 => n_654, A2 => n_650, B1 => n_652, B2 => FE_PHN80_framebuffer_buf_64_2959, ZN => n_651);
  g24893 : MOAI22D0BWP7T port map(A1 => n_654, A2 => n_648, B1 => n_652, B2 => FE_PHN104_framebuffer_buf_65_2960, ZN => n_649);
  g24894 : MOAI22D0BWP7T port map(A1 => n_645, A2 => n_653, B1 => n_644, B2 => FE_PHN161_framebuffer_buf_99_2994, ZN => n_647);
  g24896 : MOAI22D0BWP7T port map(A1 => n_645, A2 => n_648, B1 => n_644, B2 => FE_PHN183_framebuffer_buf_101_2996, ZN => n_646);
  g24895 : MOAI22D0BWP7T port map(A1 => n_645, A2 => n_650, B1 => n_644, B2 => FE_PHN26_framebuffer_buf_100_2995, ZN => n_643);
  g24897 : MOAI22D0BWP7T port map(A1 => n_645, A2 => n_641, B1 => n_644, B2 => FE_PHN113_framebuffer_buf_98_2993, ZN => n_642);
  g24886 : MOAI22D0BWP7T port map(A1 => n_659, A2 => n_641, B1 => n_658, B2 => framebuffer_buf_136_3031, ZN => n_640);
  new_counter_reg_6 : LHQD1BWP7T port map(D => n_1821, E => n_577, Q => new_counter(6));
  g24898 : MOAI22D0BWP7T port map(A1 => n_635, A2 => n_637, B1 => n_634, B2 => framebuffer_buf_128_3023, ZN => n_639);
  g24900 : MOAI22D0BWP7T port map(A1 => n_632, A2 => n_637, B1 => n_630, B2 => FE_PHN39_framebuffer_buf_54_2949, ZN => n_638);
  g24899 : MOAI22D0BWP7T port map(A1 => n_635, A2 => n_631, B1 => n_634, B2 => framebuffer_buf_129_3024, ZN => n_636);
  g24901 : MOAI22D0BWP7T port map(A1 => n_632, A2 => n_631, B1 => n_630, B2 => framebuffer_buf_55_2950, ZN => n_633);
  g24902 : MOAI22D0BWP7T port map(A1 => n_635, A2 => n_641, B1 => n_634, B2 => FE_PHN132_framebuffer_buf_124_3019, ZN => n_629);
  g24925 : MOAI22D0BWP7T port map(A1 => n_626, A2 => n_578, B1 => n_624, B2 => FE_PHN24_framebuffer_buf_61_2956, ZN => n_628);
  g24924 : MOAI22D0BWP7T port map(A1 => n_626, A2 => n_625, B1 => n_624, B2 => FE_PHN72_framebuffer_buf_60_2955, ZN => n_627);
  g24923 : MOAI22D0BWP7T port map(A1 => n_613, A2 => n_648, B1 => n_612, B2 => FE_PHN73_framebuffer_buf_151_3046, ZN => n_623);
  new_sqi_address_reg_3 : LHQD1BWP7T port map(D => n_483, E => n_681, Q => new_sqi_address(3));
  g24903 : MOAI22D0BWP7T port map(A1 => n_635, A2 => n_653, B1 => n_634, B2 => FE_PHN46_framebuffer_buf_125_3020, ZN => n_622);
  new_sqi_address_reg_8 : LHQD1BWP7T port map(D => n_460, E => n_681, Q => new_sqi_address(8));
  g24904 : MOAI22D0BWP7T port map(A1 => n_635, A2 => n_650, B1 => n_634, B2 => FE_PHN170_framebuffer_buf_126_3021, ZN => n_621);
  g24905 : MOAI22D0BWP7T port map(A1 => n_635, A2 => n_648, B1 => n_634, B2 => FE_PHN173_framebuffer_buf_127_3022, ZN => n_620);
  g24906 : MOAI22D0BWP7T port map(A1 => n_632, A2 => n_641, B1 => n_630, B2 => FE_PHN51_framebuffer_buf_50_2945, ZN => n_619);
  g24907 : MOAI22D0BWP7T port map(A1 => n_632, A2 => n_653, B1 => n_630, B2 => FE_PHN91_framebuffer_buf_51_2946, ZN => n_618);
  g24817 : MOAI22D0BWP7T port map(A1 => n_610, A2 => n_653, B1 => n_609, B2 => FE_PHN123_framebuffer_buf_111_3006, ZN => n_617);
  g24908 : MOAI22D0BWP7T port map(A1 => n_632, A2 => n_650, B1 => n_630, B2 => FE_PHN99_framebuffer_buf_52_2947, ZN => n_616);
  g24909 : MOAI22D0BWP7T port map(A1 => n_632, A2 => n_648, B1 => n_630, B2 => FE_PHN153_framebuffer_buf_53_2948, ZN => n_615);
  g24910 : MOAI22D0BWP7T port map(A1 => n_613, A2 => n_637, B1 => n_612, B2 => FE_PHN165_framebuffer_buf_152_3047, ZN => n_614);
  g24818 : MOAI22D0BWP7T port map(A1 => n_610, A2 => n_641, B1 => n_609, B2 => FE_PHN103_framebuffer_buf_110_3005, ZN => n_611);
  g24911 : MOAI22D0BWP7T port map(A1 => n_613, A2 => n_631, B1 => n_612, B2 => FE_PHN126_framebuffer_buf_153_3048, ZN => n_608);
  g24816 : MOAI22D0BWP7T port map(A1 => n_541, A2 => n_631, B1 => n_540, B2 => FE_PHN11_framebuffer_buf_91_2986, ZN => n_607);
  g24912 : MOAI22D0BWP7T port map(A1 => n_626, A2 => n_596, B1 => n_624, B2 => FE_PHN65_framebuffer_buf_56_2951, ZN => n_606);
  g24913 : MOAI22D0BWP7T port map(A1 => n_626, A2 => n_592, B1 => n_624, B2 => FE_PHN27_framebuffer_buf_57_2952, ZN => n_605);
  g24819 : MOAI22D0BWP7T port map(A1 => n_601, A2 => n_648, B1 => n_600, B2 => FE_PHN105_framebuffer_buf_77_2972, ZN => n_604);
  g24914 : MOAI22D0BWP7T port map(A1 => n_626, A2 => n_590, B1 => n_624, B2 => framebuffer_buf_58_2953, ZN => n_603);
  g24820 : MOAI22D0BWP7T port map(A1 => n_601, A2 => n_650, B1 => n_600, B2 => FE_PHN124_framebuffer_buf_76_2971, ZN => n_602);
  g24915 : MOAI22D0BWP7T port map(A1 => n_626, A2 => n_587, B1 => n_624, B2 => FE_PHN6_framebuffer_buf_59_2954, ZN => n_599);
  g24916 : MOAI22D0BWP7T port map(A1 => n_597, A2 => n_596, B1 => n_595, B2 => framebuffer_buf_130_3025, ZN => n_598);
  g24821 : MOAI22D0BWP7T port map(A1 => n_601, A2 => n_653, B1 => n_600, B2 => FE_PHN93_framebuffer_buf_75_2970, ZN => n_594);
  g24917 : MOAI22D0BWP7T port map(A1 => n_597, A2 => n_592, B1 => n_595, B2 => FE_PHN182_framebuffer_buf_131_3026, ZN => n_593);
  g24918 : MOAI22D0BWP7T port map(A1 => n_597, A2 => n_590, B1 => n_595, B2 => framebuffer_buf_132_3027, ZN => n_591);
  g24822 : MOAI22D0BWP7T port map(A1 => n_601, A2 => n_641, B1 => n_600, B2 => FE_PHN47_framebuffer_buf_74_2969, ZN => n_589);
  g24919 : MOAI22D0BWP7T port map(A1 => n_597, A2 => n_587, B1 => n_595, B2 => framebuffer_buf_133_3028, ZN => n_588);
  g24920 : MOAI22D0BWP7T port map(A1 => n_613, A2 => n_641, B1 => n_612, B2 => FE_PHN77_framebuffer_buf_148_3043, ZN => n_586);
  g24823 : MOAI22D0BWP7T port map(A1 => n_582, A2 => n_587, B1 => n_581, B2 => framebuffer_buf_157_3052, ZN => n_585);
  g24921 : MOAI22D0BWP7T port map(A1 => n_613, A2 => n_653, B1 => n_612, B2 => framebuffer_buf_149_3044, ZN => n_584);
  g24824 : MOAI22D0BWP7T port map(A1 => n_582, A2 => n_590, B1 => n_581, B2 => FE_PHN147_framebuffer_buf_156_3051, ZN => n_583);
  g24922 : MOAI22D0BWP7T port map(A1 => n_613, A2 => n_650, B1 => n_612, B2 => FE_PHN199_framebuffer_buf_150_3045, ZN => n_580);
  g24927 : MOAI22D0BWP7T port map(A1 => n_597, A2 => n_578, B1 => n_595, B2 => framebuffer_buf_135_3030, ZN => n_579);
  new_counter_reg_7 : LHQD1BWP7T port map(D => n_491, E => n_577, Q => new_counter(7));
  g24928 : MOAI22D0BWP7T port map(A1 => n_574, A2 => n_596, B1 => n_573, B2 => FE_PHN181_framebuffer_buf_104_2999, ZN => n_576);
  g24929 : MOAI22D0BWP7T port map(A1 => n_574, A2 => n_592, B1 => n_573, B2 => FE_PHN115_framebuffer_buf_105_3000, ZN => n_575);
  g24831 : OAI211D0BWP7T port map(A1 => counter(7), A2 => n_219, B => n_411, C => n_329, ZN => n_572);
  g24930 : MOAI22D0BWP7T port map(A1 => n_574, A2 => n_590, B1 => n_573, B2 => FE_PHN184_framebuffer_buf_106_3001, ZN => n_571);
  g24931 : MOAI22D0BWP7T port map(A1 => n_574, A2 => n_587, B1 => n_573, B2 => FE_PHN42_framebuffer_buf_107_3002, ZN => n_570);
  g24932 : MOAI22D0BWP7T port map(A1 => n_574, A2 => n_625, B1 => n_573, B2 => FE_PHN61_framebuffer_buf_108_3003, ZN => n_569);
  g24933 : MOAI22D0BWP7T port map(A1 => n_574, A2 => n_578, B1 => n_573, B2 => FE_PHN78_framebuffer_buf_109_3004, ZN => n_568);
  g24934 : MOAI22D0BWP7T port map(A1 => n_561, A2 => n_596, B1 => n_560, B2 => FE_PHN193_framebuffer_buf_80_2975, ZN => n_567);
  g24833 : MOAI22D0BWP7T port map(A1 => n_564, A2 => n_637, B1 => n_563, B2 => FE_PHN129_framebuffer_buf_96_2991, ZN => n_566);
  g24834 : MOAI22D0BWP7T port map(A1 => n_564, A2 => n_631, B1 => n_563, B2 => FE_PHN55_framebuffer_buf_97_2992, ZN => n_565);
  g24935 : MOAI22D0BWP7T port map(A1 => n_561, A2 => n_592, B1 => n_560, B2 => FE_PHN7_framebuffer_buf_81_2976, ZN => n_562);
  g24835 : MOAI22D0BWP7T port map(A1 => n_564, A2 => n_641, B1 => n_563, B2 => FE_PHN29_framebuffer_buf_92_2987, ZN => n_559);
  g24936 : MOAI22D0BWP7T port map(A1 => n_561, A2 => n_590, B1 => n_560, B2 => FE_PHN10_framebuffer_buf_82_2977, ZN => n_558);
  g24937 : MOAI22D0BWP7T port map(A1 => n_561, A2 => n_587, B1 => n_560, B2 => FE_PHN130_framebuffer_buf_83_2978, ZN => n_557);
  g24938 : MOAI22D0BWP7T port map(A1 => n_561, A2 => n_625, B1 => n_560, B2 => FE_PHN163_framebuffer_buf_84_2979, ZN => n_556);
  g24836 : MOAI22D0BWP7T port map(A1 => n_564, A2 => n_653, B1 => n_563, B2 => FE_PHN187_framebuffer_buf_93_2988, ZN => n_555);
  g24939 : MOAI22D0BWP7T port map(A1 => n_561, A2 => n_578, B1 => n_560, B2 => framebuffer_buf_85_2980, ZN => n_554);
  g24837 : MOAI22D0BWP7T port map(A1 => n_564, A2 => n_650, B1 => n_563, B2 => FE_PHN58_framebuffer_buf_94_2989, ZN => n_553);
  g24838 : MOAI22D0BWP7T port map(A1 => n_564, A2 => n_648, B1 => n_563, B2 => FE_PHN79_framebuffer_buf_95_2990, ZN => n_552);
  g24839 : MOAI22D0BWP7T port map(A1 => n_549, A2 => n_637, B1 => n_548, B2 => FE_PHN159_framebuffer_buf_122_3017, ZN => n_551);
  g24840 : MOAI22D0BWP7T port map(A1 => n_549, A2 => n_631, B1 => n_548, B2 => framebuffer_buf_123_3018, ZN => n_550);
  g24841 : MOAI22D0BWP7T port map(A1 => n_549, A2 => n_641, B1 => n_548, B2 => FE_PHN150_framebuffer_buf_118_3013, ZN => n_547);
  g24842 : MOAI22D0BWP7T port map(A1 => n_549, A2 => n_653, B1 => n_548, B2 => framebuffer_buf_119_3014, ZN => n_546);
  g24843 : MOAI22D0BWP7T port map(A1 => n_549, A2 => n_650, B1 => n_548, B2 => framebuffer_buf_120_3015, ZN => n_545);
  g24844 : MOAI22D0BWP7T port map(A1 => n_549, A2 => n_648, B1 => n_548, B2 => FE_PHN33_framebuffer_buf_121_3016, ZN => n_544);
  g24980 : OAI221D0BWP7T port map(A1 => n_362, A2 => n_393, B1 => n_358, B2 => n_301, C => n_486, ZN => n_543);
  g24845 : MOAI22D0BWP7T port map(A1 => n_541, A2 => n_637, B1 => n_540, B2 => FE_PHN12_framebuffer_buf_90_2985, ZN => n_542);
  g24846 : MOAI22D0BWP7T port map(A1 => n_582, A2 => n_592, B1 => n_581, B2 => framebuffer_buf_155_3050, ZN => n_539);
  g24847 : MOAI22D0BWP7T port map(A1 => n_536, A2 => n_637, B1 => n_535, B2 => FE_PHN168_framebuffer_buf_146_3041, ZN => n_538);
  g24848 : MOAI22D0BWP7T port map(A1 => n_536, A2 => n_631, B1 => n_535, B2 => FE_PHN120_framebuffer_buf_147_3042, ZN => n_537);
  g24849 : MOAI22D0BWP7T port map(A1 => n_532, A2 => n_637, B1 => n_531, B2 => FE_PHN131_framebuffer_buf_72_2967, ZN => n_534);
  g24850 : MOAI22D0BWP7T port map(A1 => n_532, A2 => n_631, B1 => n_531, B2 => FE_PHN63_framebuffer_buf_73_2968, ZN => n_533);
  g24851 : MOAI22D0BWP7T port map(A1 => n_541, A2 => n_641, B1 => n_540, B2 => FE_PHN158_framebuffer_buf_86_2981, ZN => n_530);
  g24852 : MOAI22D0BWP7T port map(A1 => n_541, A2 => n_653, B1 => n_540, B2 => FE_PHN110_framebuffer_buf_87_2982, ZN => n_529);
  g24853 : MOAI22D0BWP7T port map(A1 => n_541, A2 => n_650, B1 => n_540, B2 => FE_PHN138_framebuffer_buf_88_2983, ZN => n_528);
  g24854 : MOAI22D0BWP7T port map(A1 => n_541, A2 => n_648, B1 => n_540, B2 => FE_PHN179_framebuffer_buf_89_2984, ZN => n_527);
  g24855 : MOAI22D0BWP7T port map(A1 => n_536, A2 => n_641, B1 => n_535, B2 => FE_PHN127_framebuffer_buf_142_3037, ZN => n_526);
  g24856 : MOAI22D0BWP7T port map(A1 => n_536, A2 => n_653, B1 => n_535, B2 => FE_PHN139_framebuffer_buf_143_3038, ZN => n_525);
  g24857 : MOAI22D0BWP7T port map(A1 => n_536, A2 => n_650, B1 => n_535, B2 => FE_PHN116_framebuffer_buf_144_3039, ZN => n_524);
  g24858 : MOAI22D0BWP7T port map(A1 => n_536, A2 => n_648, B1 => n_535, B2 => FE_PHN92_framebuffer_buf_145_3040, ZN => n_523);
  g24859 : MOAI22D0BWP7T port map(A1 => n_532, A2 => n_641, B1 => n_531, B2 => FE_PHN74_framebuffer_buf_68_2963, ZN => n_522);
  g24860 : MOAI22D0BWP7T port map(A1 => n_532, A2 => n_653, B1 => n_531, B2 => FE_PHN89_framebuffer_buf_69_2964, ZN => n_521);
  g24861 : MOAI22D0BWP7T port map(A1 => n_532, A2 => n_650, B1 => n_531, B2 => FE_PHN154_framebuffer_buf_70_2965, ZN => n_520);
  g24862 : MOAI22D0BWP7T port map(A1 => n_532, A2 => n_648, B1 => n_531, B2 => framebuffer_buf_71_2966, ZN => n_519);
  g24863 : MOAI22D0BWP7T port map(A1 => n_601, A2 => n_637, B1 => n_600, B2 => FE_PHN142_framebuffer_buf_78_2973, ZN => n_518);
  g24864 : MOAI22D0BWP7T port map(A1 => n_601, A2 => n_631, B1 => n_600, B2 => FE_PHN157_framebuffer_buf_79_2974, ZN => n_517);
  g24865 : MOAI22D0BWP7T port map(A1 => n_610, A2 => n_637, B1 => n_609, B2 => FE_PHN118_framebuffer_buf_114_3009, ZN => n_516);
  g24866 : MOAI22D0BWP7T port map(A1 => n_610, A2 => n_631, B1 => n_609, B2 => framebuffer_buf_115_3010, ZN => n_515);
  g24867 : MOAI22D0BWP7T port map(A1 => n_582, A2 => n_596, B1 => n_581, B2 => FE_PHN190_framebuffer_buf_154_3049, ZN => n_514);
  g24878 : MOAI22D0BWP7T port map(A1 => n_610, A2 => n_650, B1 => n_609, B2 => FE_PHN122_framebuffer_buf_112_3007, ZN => n_513);
  g24879 : MOAI22D0BWP7T port map(A1 => n_610, A2 => n_648, B1 => n_609, B2 => framebuffer_buf_113_3008, ZN => n_512);
  g24880 : MOAI22D0BWP7T port map(A1 => n_659, A2 => n_637, B1 => n_658, B2 => FE_PHN81_framebuffer_buf_140_3035, ZN => n_511);
  g24881 : MOAI22D0BWP7T port map(A1 => n_659, A2 => n_631, B1 => n_658, B2 => FE_PHN102_framebuffer_buf_141_3036, ZN => n_510);
  g24882 : MOAI22D0BWP7T port map(A1 => n_654, A2 => n_637, B1 => n_652, B2 => FE_PHN48_framebuffer_buf_66_2961, ZN => n_509);
  g24883 : MOAI22D0BWP7T port map(A1 => n_654, A2 => n_631, B1 => n_652, B2 => FE_PHN107_framebuffer_buf_67_2962, ZN => n_508);
  g24884 : MOAI22D0BWP7T port map(A1 => n_645, A2 => n_637, B1 => n_644, B2 => FE_PHN60_framebuffer_buf_102_2997, ZN => n_507);
  g24885 : MOAI22D0BWP7T port map(A1 => n_645, A2 => n_631, B1 => n_644, B2 => FE_PHN156_framebuffer_buf_103_2998, ZN => n_506);
  g25071 : OAI211D0BWP7T port map(A1 => n_504, A2 => n_181, B => n_376, C => n_207, ZN => n_505);
  g25030 : AOI211D0BWP7T port map(A1 => n_375, A2 => n_26, B => n_378, C => n_356, ZN => n_503);
  g24779 : MOAI22D0BWP7T port map(A1 => n_500, A2 => n_650, B1 => n_499, B2 => FE_PHN30_calc_buf_out_4_2875, ZN => n_502);
  g24780 : MOAI22D0BWP7T port map(A1 => n_500, A2 => n_653, B1 => n_499, B2 => FE_PHN28_calc_buf_out_3_2874, ZN => n_501);
  g24781 : MOAI22D0BWP7T port map(A1 => n_500, A2 => n_641, B1 => n_499, B2 => FE_PHN188_calc_buf_out_2_2873, ZN => n_498);
  g24782 : MOAI22D0BWP7T port map(A1 => n_500, A2 => n_631, B1 => n_499, B2 => FE_PHN84_calc_buf_out_7_2878, ZN => n_497);
  g24783 : MOAI22D0BWP7T port map(A1 => n_500, A2 => n_637, B1 => n_499, B2 => FE_PHN83_calc_buf_out_6_2877, ZN => n_496);
  g24786 : AO22D0BWP7T port map(A1 => n_499, A2 => FE_PHN14_calc_buf_out_1_2872, B1 => sqi_data_in(1), B2 => n_493, Z => n_495);
  g24787 : AO22D0BWP7T port map(A1 => n_499, A2 => FE_PHN13_calc_buf_out_0_2871, B1 => sqi_data_in(0), B2 => n_493, Z => n_494);
  g24778 : MOAI22D0BWP7T port map(A1 => n_500, A2 => n_648, B1 => n_499, B2 => FE_PHN37_calc_buf_out_5_2876, ZN => n_492);
  g24981 : OAI32D0BWP7T port map(A1 => counter(7), A2 => n_324, A3 => n_380, B1 => n_504, B2 => n_326, ZN => n_491);
  new_sqi_address_reg_0 : LHQD1BWP7T port map(D => n_350, E => n_681, Q => new_sqi_address(0));
  g25012 : MOAI22D0BWP7T port map(A1 => n_477, A2 => n_637, B1 => n_476, B2 => FE_PHN100_framebuffer_buf_42_2937, ZN => n_490);
  new_sqi_address_reg_5 : LHQD1BWP7T port map(D => n_333, E => n_681, Q => new_sqi_address(5));
  new_sqi_address_reg_2 : LHQD1BWP7T port map(D => n_396, E => n_681, Q => new_sqi_address(2));
  g25096 : AOI221D0BWP7T port map(A1 => n_488, A2 => sqi_address(9), B1 => n_459, B2 => n_32, C => n_310, ZN => n_489);
  g25098 : AOI221D0BWP7T port map(A1 => n_158, A2 => n_237, B1 => n_361, B2 => n_410, C => n_308, ZN => n_486);
  g25099 : NR3D0BWP7T port map(A1 => n_364, A2 => n_315, A3 => n_259, ZN => n_485);
  g25143 : OAI211D0BWP7T port map(A1 => n_242, A2 => n_262, B => n_306, C => n_419, ZN => n_484);
  g24940 : OAI211D0BWP7T port map(A1 => n_204, A2 => n_106, B => n_323, C => n_215, ZN => n_483);
  g24964 : INVD5BWP7T port map(I => n_700, ZN => single);
  g24966 : INVD5BWP7T port map(I => n_699, ZN => sqi_rw);
  new_counter_reg_5 : LHQD1BWP7T port map(D => n_381, E => n_577, Q => new_counter(5));
  g25011 : MOAI22D0BWP7T port map(A1 => n_470, A2 => n_648, B1 => n_469, B2 => framebuffer_buf_23_2918, ZN => n_479);
  g24996 : MOAI22D0BWP7T port map(A1 => n_477, A2 => n_648, B1 => n_476, B2 => framebuffer_buf_41_2936, ZN => n_478);
  g25000 : MOAI22D0BWP7T port map(A1 => n_473, A2 => n_637, B1 => n_472, B2 => FE_PHN88_framebuffer_buf_48_2943, ZN => n_475);
  g25001 : MOAI22D0BWP7T port map(A1 => n_473, A2 => n_631, B1 => n_472, B2 => FE_PHN149_framebuffer_buf_49_2944, ZN => n_474);
  g25002 : MOAI22D0BWP7T port map(A1 => n_470, A2 => n_637, B1 => n_469, B2 => FE_PHN185_framebuffer_buf_24_2919, ZN => n_471);
  g25003 : MOAI22D0BWP7T port map(A1 => n_470, A2 => n_631, B1 => n_469, B2 => FE_PHN86_framebuffer_buf_25_2920, ZN => n_468);
  g25004 : MOAI22D0BWP7T port map(A1 => n_473, A2 => n_641, B1 => n_472, B2 => FE_PHN144_framebuffer_buf_44_2939, ZN => n_467);
  g25005 : MOAI22D0BWP7T port map(A1 => n_473, A2 => n_653, B1 => n_472, B2 => FE_PHN52_framebuffer_buf_45_2940, ZN => n_466);
  g25006 : MOAI22D0BWP7T port map(A1 => n_473, A2 => n_650, B1 => n_472, B2 => FE_PHN106_framebuffer_buf_46_2941, ZN => n_465);
  g25007 : MOAI22D0BWP7T port map(A1 => n_473, A2 => n_648, B1 => n_472, B2 => FE_PHN145_framebuffer_buf_47_2942, ZN => n_464);
  g25008 : MOAI22D0BWP7T port map(A1 => n_470, A2 => n_641, B1 => n_469, B2 => FE_PHN18_framebuffer_buf_20_2915, ZN => n_463);
  g25009 : MOAI22D0BWP7T port map(A1 => n_470, A2 => n_653, B1 => n_469, B2 => FE_PHN67_framebuffer_buf_21_2916, ZN => n_462);
  g25010 : MOAI22D0BWP7T port map(A1 => n_470, A2 => n_650, B1 => n_469, B2 => FE_PHN76_framebuffer_buf_22_2917, ZN => n_461);
  g25049 : AO221D0BWP7T port map(A1 => n_459, A2 => n_41, B1 => n_488, B2 => sqi_address(8), C => n_374, Z => n_460);
  g25014 : MOAI22D0BWP7T port map(A1 => n_455, A2 => n_637, B1 => n_454, B2 => FE_PHN82_framebuffer_buf_18_2913, ZN => n_457);
  g25015 : MOAI22D0BWP7T port map(A1 => n_455, A2 => n_631, B1 => n_454, B2 => FE_PHN95_framebuffer_buf_19_2914, ZN => n_456);
  g25016 : MOAI22D0BWP7T port map(A1 => n_477, A2 => n_641, B1 => n_476, B2 => FE_PHN35_framebuffer_buf_38_2933, ZN => n_453);
  g25017 : MOAI22D0BWP7T port map(A1 => n_477, A2 => n_653, B1 => n_476, B2 => FE_PHN96_framebuffer_buf_39_2934, ZN => n_452);
  g25018 : MOAI22D0BWP7T port map(A1 => n_477, A2 => n_650, B1 => n_476, B2 => FE_PHN160_framebuffer_buf_40_2935, ZN => n_451);
  g25020 : MOAI22D0BWP7T port map(A1 => n_455, A2 => n_641, B1 => n_454, B2 => FE_PHN133_framebuffer_buf_14_2909, ZN => n_450);
  g25021 : MOAI22D0BWP7T port map(A1 => n_455, A2 => n_653, B1 => n_454, B2 => FE_PHN98_framebuffer_buf_15_2910, ZN => n_449);
  g25022 : MOAI22D0BWP7T port map(A1 => n_455, A2 => n_650, B1 => n_454, B2 => FE_PHN85_framebuffer_buf_16_2911, ZN => n_448);
  g25023 : MOAI22D0BWP7T port map(A1 => n_455, A2 => n_648, B1 => n_454, B2 => framebuffer_buf_17_2912, ZN => n_447);
  g25024 : MOAI22D0BWP7T port map(A1 => n_444, A2 => n_637, B1 => n_443, B2 => FE_PHN22_framebuffer_buf_30_2925, ZN => n_446);
  g25025 : MOAI22D0BWP7T port map(A1 => n_444, A2 => n_631, B1 => n_443, B2 => FE_PHN44_framebuffer_buf_31_2926, ZN => n_445);
  g25026 : MOAI22D0BWP7T port map(A1 => n_444, A2 => n_641, B1 => n_443, B2 => FE_PHN41_framebuffer_buf_26_2921, ZN => n_442);
  g25027 : MOAI22D0BWP7T port map(A1 => n_444, A2 => n_653, B1 => n_443, B2 => FE_PHN117_framebuffer_buf_27_2922, ZN => n_441);
  g25028 : MOAI22D0BWP7T port map(A1 => n_444, A2 => n_650, B1 => n_443, B2 => framebuffer_buf_28_2923, ZN => n_440);
  g25029 : MOAI22D0BWP7T port map(A1 => n_444, A2 => n_648, B1 => n_443, B2 => FE_PHN20_framebuffer_buf_29_2924, ZN => n_439);
  g25031 : MOAI22D0BWP7T port map(A1 => n_436, A2 => n_592, B1 => n_435, B2 => FE_PHN45_framebuffer_buf_9_2904, ZN => n_438);
  g25032 : MOAI22D0BWP7T port map(A1 => n_436, A2 => n_590, B1 => n_435, B2 => FE_PHN38_framebuffer_buf_10_2905, ZN => n_437);
  g25033 : MOAI22D0BWP7T port map(A1 => n_436, A2 => n_587, B1 => n_435, B2 => FE_PHN53_framebuffer_buf_11_2906, ZN => n_434);
  g25034 : MOAI22D0BWP7T port map(A1 => n_436, A2 => n_625, B1 => n_435, B2 => FE_PHN136_framebuffer_buf_12_2907, ZN => n_433);
  g25035 : MOAI22D0BWP7T port map(A1 => n_436, A2 => n_578, B1 => n_435, B2 => FE_PHN134_framebuffer_buf_13_2908, ZN => n_432);
  g25036 : MOAI22D0BWP7T port map(A1 => n_429, A2 => n_596, B1 => n_428, B2 => FE_PHN34_framebuffer_buf_32_2927, ZN => n_431);
  g25037 : MOAI22D0BWP7T port map(A1 => n_429, A2 => n_592, B1 => n_428, B2 => FE_PHN112_framebuffer_buf_33_2928, ZN => n_430);
  g25038 : MOAI22D0BWP7T port map(A1 => n_429, A2 => n_590, B1 => n_428, B2 => FE_PHN90_framebuffer_buf_34_2929, ZN => n_427);
  g25039 : MOAI22D0BWP7T port map(A1 => n_429, A2 => n_587, B1 => n_428, B2 => FE_PHN57_framebuffer_buf_35_2930, ZN => n_426);
  g25040 : MOAI22D0BWP7T port map(A1 => n_429, A2 => n_625, B1 => n_428, B2 => FE_PHN70_framebuffer_buf_36_2931, ZN => n_425);
  g25041 : MOAI22D0BWP7T port map(A1 => n_429, A2 => n_578, B1 => n_428, B2 => framebuffer_buf_37_2932, ZN => n_424);
  g25042 : MOAI22D0BWP7T port map(A1 => n_436, A2 => n_596, B1 => n_435, B2 => FE_PHN101_framebuffer_buf_8_2903, ZN => n_423);
  g25047 : AOI222D0BWP7T port map(A1 => n_360, A2 => counter(5), B1 => n_409, B2 => n_38, C1 => n_193, C2 => counter(3), ZN => n_422);
  g25013 : MOAI22D0BWP7T port map(A1 => n_477, A2 => n_631, B1 => n_476, B2 => FE_PHN140_framebuffer_buf_43_2938, ZN => n_421);
  g25110 : OAI221D0BWP7T port map(A1 => n_419, A2 => n_234, B1 => n_418, B2 => n_371, C => n_261, ZN => n_420);
  g24954 : INVD5BWP7T port map(I => n_702, ZN => sqi_data_out(1));
  g24952 : INVD5BWP7T port map(I => n_703, ZN => sqi_data_out(2));
  g24950 : INVD5BWP7T port map(I => n_704, ZN => sqi_data_out(4));
  g24948 : INVD5BWP7T port map(I => n_705, ZN => sqi_data_out(3));
  g24946 : INVD5BWP7T port map(I => n_706, ZN => sqi_data_out(6));
  new_sqi_address_reg_7 : LHQD1BWP7T port map(D => n_305, E => n_681, Q => new_sqi_address(7));
  g24944 : INVD5BWP7T port map(I => n_707, ZN => sqi_data_out(5));
  g25085 : AOI33D0BWP7T port map(A1 => n_263, A2 => n_410, A3 => n_504, B1 => n_409, B2 => n_75, B3 => counter(7), ZN => n_411);
  g25134 : AOI221D0BWP7T port map(A1 => n_366, A2 => n_410, B1 => n_488, B2 => sqi_address(14), C => n_265, ZN => n_408);
  new_sqi_address_reg_1 : LHQD1BWP7T port map(D => n_313, E => n_681, Q => new_sqi_address(1));
  g25136 : ND2D0BWP7T port map(A1 => n_303, A2 => n_504, ZN => n_674);
  g25062 : ND2D1BWP7T port map(A1 => n_406, A2 => n_401, ZN => n_540);
  g25063 : ND2D1BWP7T port map(A1 => n_406, A2 => n_405, ZN => n_560);
  g25067 : ND2D1BWP7T port map(A1 => n_404, A2 => n_405, ZN => n_624);
  g25066 : ND2D1BWP7T port map(A1 => n_404, A2 => n_403, ZN => n_630);
  g25065 : ND2D1BWP7T port map(A1 => n_398, A2 => n_403, ZN => n_644);
  g25064 : ND2D1BWP7T port map(A1 => n_406, A2 => n_400, ZN => n_563);
  new_counter_reg_3 : LHQD1BWP7T port map(D => n_328, E => n_577, Q => new_counter(3));
  single_reg : LHD1BWP7T port map(D => n_54, E => n_402, Q => UNCONNECTED, QN => n_700);
  sqi_rw_reg : LHD1BWP7T port map(D => n_138, E => n_402, Q => UNCONNECTED0, QN => n_699);
  new_counter_reg_2 : LHQD1BWP7T port map(D => n_281, E => n_577, Q => new_counter(2));
  new_counter_reg_0 : LHQD1BWP7T port map(D => n_253, E => n_577, Q => new_counter(0));
  new_counter_reg_4 : LHQD1BWP7T port map(D => n_284, E => n_577, Q => new_counter(4));
  new_counter_reg_1 : LHQD1BWP7T port map(D => n_248, E => n_577, Q => new_counter(1));
  g25050 : ND2D1BWP7T port map(A1 => n_399, A2 => n_405, ZN => n_581);
  g25051 : ND2D1BWP7T port map(A1 => n_404, A2 => n_401, ZN => n_652);
  g25052 : ND2D1BWP7T port map(A1 => n_404, A2 => n_400, ZN => n_531);
  g25053 : ND2D1BWP7T port map(A1 => n_399, A2 => n_403, ZN => n_612);
  g25054 : ND2D1BWP7T port map(A1 => n_398, A2 => n_401, ZN => n_609);
  g25055 : ND2D1BWP7T port map(A1 => n_406, A2 => n_403, ZN => n_600);
  g25056 : ND2D1BWP7T port map(A1 => n_397, A2 => n_403, ZN => n_634);
  g25057 : ND2D1BWP7T port map(A1 => n_397, A2 => n_405, ZN => n_595);
  g25058 : ND2D1BWP7T port map(A1 => n_397, A2 => n_401, ZN => n_658);
  g25059 : ND2D1BWP7T port map(A1 => n_397, A2 => n_400, ZN => n_535);
  g25060 : ND2D1BWP7T port map(A1 => n_398, A2 => n_405, ZN => n_573);
  g25061 : ND2D1BWP7T port map(A1 => n_398, A2 => n_400, ZN => n_548);
  new_sqi_address_reg_6 : LHQD1BWP7T port map(D => n_274, E => n_681, Q => new_sqi_address(6));
  g25074 : AO221D0BWP7T port map(A1 => n_213, A2 => y(2), B1 => n_488, B2 => sqi_address(2), C => n_278, Z => n_396);
  g25081 : MOAI22D0BWP7T port map(A1 => n_386, A2 => n_648, B1 => n_390, B2 => FE_PHN166_framebuffer_buf_5_2900, ZN => n_392);
  g25083 : AO22D0BWP7T port map(A1 => n_390, A2 => FE_PHN40_framebuffer_buf_0_2895, B1 => sqi_data_in(0), B2 => n_388, Z => n_391);
  g25084 : AO22D0BWP7T port map(A1 => n_390, A2 => FE_PHN43_framebuffer_buf_1_2896, B1 => sqi_data_in(1), B2 => n_388, Z => n_389);
  g25086 : MOAI22D0BWP7T port map(A1 => n_386, A2 => n_637, B1 => n_390, B2 => FE_PHN111_framebuffer_buf_6_2901, ZN => n_387);
  g25087 : MOAI22D0BWP7T port map(A1 => n_386, A2 => n_631, B1 => n_390, B2 => FE_PHN9_framebuffer_buf_7_2902, ZN => n_385);
  g25088 : MOAI22D0BWP7T port map(A1 => n_386, A2 => n_641, B1 => n_390, B2 => FE_PHN21_framebuffer_buf_2_2897, ZN => n_384);
  g25089 : MOAI22D0BWP7T port map(A1 => n_386, A2 => n_653, B1 => n_390, B2 => framebuffer_buf_3_2898, ZN => n_383);
  g25090 : MOAI22D0BWP7T port map(A1 => n_386, A2 => n_650, B1 => n_390, B2 => FE_PHN178_framebuffer_buf_4_2899, ZN => n_382);
  new_sqi_address_reg_4 : LHQD1BWP7T port map(D => n_289, E => n_681, Q => new_sqi_address(4));
  g25072 : MOAI22D0BWP7T port map(A1 => n_380, A2 => counter(5), B1 => n_379, B2 => counter(5), ZN => n_381);
  g25111 : OAI221D0BWP7T port map(A1 => n_191, A2 => n_252, B1 => n_40, B2 => n_377, C => n_186, ZN => n_378);
  g25116 : AOI31D0BWP7T port map(A1 => n_375, A2 => n_504, A3 => counter(6), B => n_276, ZN => n_376);
  g25117 : OAI32D0BWP7T port map(A1 => counter(2), A2 => n_311, A3 => n_35, B1 => n_355, B2 => n_233, ZN => n_374);
  g25127 : OAI211D0BWP7T port map(A1 => n_307, A2 => n_208, B => n_372, C => n_371, ZN => n_373);
  g25129 : OAI31D0BWP7T port map(A1 => n_309, A2 => n_369, A3 => n_264, B => n_368, ZN => n_370);
  g25139 : OA21D0BWP7T port map(A1 => n_231, A2 => n_366, B => n_410, Z => n_367);
  g25140 : AO22D0BWP7T port map(A1 => n_364, A2 => n_271, B1 => n_363, B2 => n_229, Z => n_365);
  g25145 : AOI21D0BWP7T port map(A1 => n_361, A2 => n_418, B => n_360, ZN => n_362);
  sqi_data_out_reg_6 : LND1BWP7T port map(D => n_290, EN => n_359, Q => UNCONNECTED1, QN => n_706);
  sqi_data_out_reg_5 : LND1BWP7T port map(D => n_275, EN => n_359, Q => UNCONNECTED2, QN => n_707);
  g25179 : OR2D1BWP7T port map(A1 => n_626, A2 => n_255, Z => n_654);
  g25170 : OR2D1BWP7T port map(A1 => n_626, A2 => n_358, Z => n_532);
  g24986 : AO22D0BWP7T port map(A1 => n_353, A2 => FE_PHN17_calc_buf_out_17_2888, B1 => sqi_data_in(1), B2 => n_343, Z => n_357);
  sqi_data_out_reg_4 : LND1BWP7T port map(D => n_291, EN => n_359, Q => UNCONNECTED3, QN => n_704);
  g25197 : OAI31D0BWP7T port map(A1 => n_355, A2 => n_245, A3 => n_314, B => n_267, ZN => n_356);
  sqi_data_out_reg_2 : LND1BWP7T port map(D => n_296, EN => n_359, Q => UNCONNECTED4, QN => n_703);
  sqi_data_out_reg_1 : LND1BWP7T port map(D => n_297, EN => n_359, Q => UNCONNECTED5, QN => n_702);
  g24973 : MOAI22D0BWP7T port map(A1 => n_338, A2 => n_641, B1 => n_353, B2 => FE_PHN135_calc_buf_out_18_2889, ZN => n_354);
  g24975 : ND4D0BWP7T port map(A1 => n_241, A2 => n_136, A3 => n_320, A4 => FE_OFN2_n_0, ZN => n_352);
  g24977 : MOAI22D0BWP7T port map(A1 => n_341, A2 => n_648, B1 => n_347, B2 => FE_PHN164_calc_buf_out_13_2884, ZN => n_351);
  g24982 : AO221D0BWP7T port map(A1 => n_128, A2 => y(0), B1 => n_488, B2 => sqi_address(0), C => n_298, Z => n_350);
  g24983 : AO22D0BWP7T port map(A1 => n_347, A2 => FE_PHN186_calc_buf_out_8_2879, B1 => sqi_data_in(0), B2 => n_345, Z => n_348);
  g24984 : AO22D0BWP7T port map(A1 => n_347, A2 => calc_buf_out_9_2880, B1 => sqi_data_in(1), B2 => n_345, Z => n_346);
  g24985 : AO22D0BWP7T port map(A1 => n_353, A2 => FE_PHN15_calc_buf_out_16_2887, B1 => sqi_data_in(0), B2 => n_343, Z => n_344);
  sqi_data_out_reg_3 : LND1BWP7T port map(D => n_292, EN => n_359, Q => UNCONNECTED6, QN => n_705);
  g24987 : MOAI22D0BWP7T port map(A1 => n_341, A2 => n_637, B1 => n_347, B2 => FE_PHN75_calc_buf_out_14_2885, ZN => n_342);
  g24988 : MOAI22D0BWP7T port map(A1 => n_341, A2 => n_631, B1 => n_347, B2 => FE_PHN64_calc_buf_out_15_2886, ZN => n_340);
  g24989 : MOAI22D0BWP7T port map(A1 => n_338, A2 => n_637, B1 => n_353, B2 => FE_PHN31_calc_buf_out_22_2893, ZN => n_339);
  g24990 : MOAI22D0BWP7T port map(A1 => n_338, A2 => n_631, B1 => n_353, B2 => FE_PHN23_calc_buf_out_23_2894, ZN => n_337);
  g24991 : MOAI22D0BWP7T port map(A1 => n_341, A2 => n_641, B1 => n_347, B2 => calc_buf_out_10_2881, ZN => n_336);
  g24992 : MOAI22D0BWP7T port map(A1 => n_341, A2 => n_653, B1 => n_347, B2 => FE_PHN49_calc_buf_out_11_2882, ZN => n_335);
  g24993 : MOAI22D0BWP7T port map(A1 => n_341, A2 => n_650, B1 => n_347, B2 => FE_PHN32_calc_buf_out_12_2883, ZN => n_334);
  g25045 : ND2D0BWP7T port map(A1 => n_283, A2 => n_133, ZN => n_333);
  g24997 : MOAI22D0BWP7T port map(A1 => n_338, A2 => n_650, B1 => n_353, B2 => FE_PHN25_calc_buf_out_20_2891, ZN => n_332);
  g24998 : MOAI22D0BWP7T port map(A1 => n_338, A2 => n_648, B1 => n_353, B2 => FE_PHN152_calc_buf_out_21_2892, ZN => n_331);
  g25019 : MOAI22D0BWP7T port map(A1 => n_338, A2 => n_653, B1 => n_353, B2 => FE_PHN94_calc_buf_out_19_2890, ZN => n_330);
  g24994 : ND3D0BWP7T port map(A1 => n_285, A2 => n_109, A3 => n_15, ZN => n_499);
  g25112 : AOI22D0BWP7T port map(A1 => n_169, A2 => n_225, B1 => n_173, B2 => counter(7), ZN => n_329);
  g25073 : OAI222D0BWP7T port map(A1 => n_358, A2 => n_167, B1 => n_279, B2 => n_327, C1 => n_321, C2 => n_244, ZN => n_328);
  g25095 : AOI21D0BWP7T port map(A1 => n_325, A2 => n_324, B => n_379, ZN => n_326);
  g25118 : AOI22D0BWP7T port map(A1 => n_214, A2 => y(3), B1 => n_488, B2 => sqi_address(3), ZN => n_323);
  g25122 : AOI21D0BWP7T port map(A1 => n_321, A2 => n_319, B => n_318, ZN => n_399);
  g25091 : ND4D0BWP7T port map(A1 => n_200, A2 => n_29, A3 => n_320, A4 => n_10, ZN => n_402);
  g25123 : AOI21D0BWP7T port map(A1 => n_156, A2 => n_319, B => n_318, ZN => n_397);
  g25103 : ND2D1BWP7T port map(A1 => n_316, A2 => n_401, ZN => n_454);
  g25104 : ND2D1BWP7T port map(A1 => n_317, A2 => n_400, ZN => n_472);
  g25105 : ND2D1BWP7T port map(A1 => n_317, A2 => n_405, ZN => n_428);
  g25106 : ND2D1BWP7T port map(A1 => n_317, A2 => n_401, ZN => n_476);
  g25100 : ND2D1BWP7T port map(A1 => n_316, A2 => n_405, ZN => n_435);
  g25101 : ND2D1BWP7T port map(A1 => n_316, A2 => n_400, ZN => n_469);
  g25102 : ND2D1BWP7T port map(A1 => n_317, A2 => n_403, ZN => n_443);
  g25092 : IND4D0BWP7T port map(A1 => n_250, B1 => n_320, B2 => n_137, B3 => n_196, ZN => n_577);
  g25189 : OAI31D0BWP7T port map(A1 => counter(3), A2 => n_418, A3 => n_314, B => n_235, ZN => n_315);
  g25043 : ND3D0BWP7T port map(A1 => n_221, A2 => n_277, A3 => n_37, ZN => n_313);
  g24976 : ND4D0BWP7T port map(A1 => n_224, A2 => n_286, A3 => n_144, A4 => n_311, ZN => n_312);
  g25141 : MOAI22D0BWP7T port map(A1 => n_176, A2 => n_309, B1 => n_91, B2 => n_175, ZN => n_310);
  g25142 : OAI33D0BWP7T port map(A1 => n_309, A2 => n_80, A3 => n_302, B1 => n_393, B2 => n_307, B3 => n_311, ZN => n_308);
  g25159 : ND2D0BWP7T port map(A1 => n_364, A2 => n_393, ZN => n_306);
  g24974 : ND4D0BWP7T port map(A1 => n_205, A2 => n_212, A3 => n_97, A4 => n_148, ZN => n_305);
  g24956 : INVD5BWP7T port map(I => n_701, ZN => sqi_data_out(0));
  g25194 : OAI21D0BWP7T port map(A1 => n_302, A2 => n_57, B => n_301, ZN => n_303);
  g24942 : INVD5BWP7T port map(I => n_708, ZN => sqi_data_out(7));
  g25124 : AOI21D0BWP7T port map(A1 => n_319, A2 => counter(2), B => n_299, ZN => n_404);
  g25125 : AOI21D0BWP7T port map(A1 => n_309, A2 => n_319, B => n_318, ZN => n_398);
  g25126 : AOI21D0BWP7T port map(A1 => n_319, A2 => n_355, B => n_299, ZN => n_406);
  g25177 : ND2D1BWP7T port map(A1 => n_254, A2 => n_268, ZN => n_632);
  g25097 : NR3D0BWP7T port map(A1 => n_217, A2 => n_273, A3 => y(0), ZN => n_298);
  g25077 : AO222D0BWP7T port map(A1 => n_295, A2 => calc_buf_in(0), B1 => n_294, B2 => edit_buf_in(1), C1 => n_293, C2 => row_buf(1), Z => n_297);
  g25078 : AO222D0BWP7T port map(A1 => n_295, A2 => calc_buf_in(1), B1 => n_294, B2 => edit_buf_in(2), C1 => n_293, C2 => row_buf(2), Z => n_296);
  g25079 : AO222D0BWP7T port map(A1 => n_295, A2 => calc_buf_in(2), B1 => n_294, B2 => edit_buf_in(3), C1 => n_293, C2 => row_buf(3), Z => n_292);
  g25080 : AO222D0BWP7T port map(A1 => n_295, A2 => calc_buf_in(3), B1 => n_294, B2 => edit_buf_in(4), C1 => n_293, C2 => row_buf(4), Z => n_291);
  g25082 : AO222D0BWP7T port map(A1 => n_295, A2 => calc_buf_in(5), B1 => n_294, B2 => edit_buf_in(6), C1 => n_293, C2 => calc_buf_in(0), Z => n_290);
  g25094 : AO221D0BWP7T port map(A1 => n_163, A2 => y(4), B1 => n_488, B2 => sqi_address(4), C => n_216, Z => n_289);
  g25069 : ND3D0BWP7T port map(A1 => n_222, A2 => n_223, A3 => n_286, ZN => n_287);
  g25113 : AOI211XD0BWP7T port map(A1 => n_160, A2 => state(3), B => n_166, C => n_12, ZN => n_285);
  g25114 : OAI32D0BWP7T port map(A1 => n_240, A2 => n_227, A3 => n_280, B1 => n_70, B2 => n_238, ZN => n_284);
  g25115 : AOI22D0BWP7T port map(A1 => n_165, A2 => y(5), B1 => n_488, B2 => sqi_address(5), ZN => n_283);
  g25121 : OAI32D0BWP7T port map(A1 => counter(2), A2 => n_358, A3 => n_280, B1 => n_355, B2 => n_279, ZN => n_281);
  g25133 : NR2D0BWP7T port map(A1 => n_277, A2 => y(2), ZN => n_278);
  g25144 : OAI31D0BWP7T port map(A1 => n_324, A2 => n_363, A3 => n_116, B => n_226, ZN => n_276);
  g25068 : AO222D0BWP7T port map(A1 => n_295, A2 => calc_buf_in(4), B1 => n_294, B2 => edit_buf_in(5), C1 => n_293, C2 => row_buf(5), Z => n_275);
  g25167 : ND2D0BWP7T port map(A1 => n_174, A2 => counter(6), ZN => n_368);
  g25048 : OAI221D0BWP7T port map(A1 => n_135, A2 => n_273, B1 => n_211, B2 => n_151, C => n_95, ZN => n_274);
  g25261 : AO22D0BWP7T port map(A1 => n_375, A2 => n_393, B1 => n_271, B2 => n_269, Z => n_272);
  g25258 : MAOI22D0BWP7T port map(A1 => n_269, A2 => n_268, B1 => n_256, B2 => counter(0), ZN => n_270);
  g25221 : AOI21D0BWP7T port map(A1 => n_488, A2 => sqi_address(10), B => n_194, ZN => n_267);
  g25188 : OAI22D0BWP7T port map(A1 => n_230, A2 => n_99, B1 => n_264, B2 => n_115, ZN => n_265);
  g25193 : OAI21D0BWP7T port map(A1 => n_257, A2 => n_268, B => n_262, ZN => n_263);
  sqi_data_out_reg_7 : LND1BWP7T port map(D => n_199, EN => n_359, Q => UNCONNECTED7, QN => n_708);
  sqi_data_out_reg_0 : LND1BWP7T port map(D => n_218, EN => n_359, Q => UNCONNECTED8, QN => n_701);
  g25201 : MAOI22D0BWP7T port map(A1 => n_488, A2 => sqi_address(12), B1 => n_262, B2 => n_324, ZN => n_261);
  g25207 : OAI32D0BWP7T port map(A1 => n_309, A2 => n_358, A3 => n_311, B1 => n_258, B2 => n_257, ZN => n_259);
  g25214 : OAI22D0BWP7T port map(A1 => n_262, A2 => n_246, B1 => n_256, B2 => n_258, ZN => n_360);
  g25181 : OR2D1BWP7T port map(A1 => n_597, A2 => n_255, Z => n_659);
  g25175 : OR2D1BWP7T port map(A1 => n_561, A2 => n_255, Z => n_541);
  g25171 : OR2D1BWP7T port map(A1 => n_597, A2 => n_358, Z => n_536);
  g25173 : OR2D1BWP7T port map(A1 => n_561, A2 => n_258, Z => n_601);
  g25218 : INVD1BWP7T port map(I => n_254, ZN => n_626);
  g25076 : OAI222D0BWP7T port map(A1 => n_107, A2 => counter(1), B1 => n_252, B2 => n_247, C1 => counter(0), C2 => n_280, ZN => n_253);
  g25070 : IND4D0BWP7T port map(A1 => n_250, B1 => FE_OFN2_n_0, B2 => n_79, B3 => n_739, ZN => n_251);
  g25119 : OAI222D0BWP7T port map(A1 => n_247, A2 => n_246, B1 => n_245, B2 => n_280, C1 => n_255, C2 => n_244, ZN => n_248);
  g25128 : NR2D0BWP7T port map(A1 => n_380, A2 => n_242, ZN => n_243);
  g25131 : AOI211XD0BWP7T port map(A1 => n_121, A2 => n_111, B => n_153, C => n_11, ZN => n_241);
  g25147 : IOA21D1BWP7T port map(A1 => n_240, A2 => n_319, B => n_239, ZN => n_299);
  g25148 : OA21D0BWP7T port map(A1 => n_120, A2 => state(3), B => n_239, Z => n_316);
  g25138 : OAI21D0BWP7T port map(A1 => state(3), A2 => counter(4), B => n_239, ZN => n_318);
  g25137 : OAI21D0BWP7T port map(A1 => n_244, A2 => counter(4), B => n_238, ZN => n_379);
  g25149 : OA21D0BWP7T port map(A1 => n_237, A2 => state(3), B => n_239, Z => n_317);
  g25150 : OAI21D0BWP7T port map(A1 => n_122, A2 => state(3), B => n_239, ZN => n_390);
  g25107 : IND2D1BWP7T port map(A1 => n_236, B1 => n_405, ZN => n_347);
  g25108 : IND2D1BWP7T port map(A1 => n_236, B1 => n_401, ZN => n_353);
  g25109 : ND4D1BWP7T port map(A1 => n_146, A2 => n_102, A3 => n_319, A4 => state(2), ZN => n_681);
  g25260 : OA22D0BWP7T port map(A1 => n_155, A2 => n_234, B1 => n_255, B2 => n_256, Z => n_235);
  g25164 : OA221D0BWP7T port map(A1 => n_203, A2 => n_246, B1 => counter(0), B2 => n_147, C => n_232, Z => n_233);
  g25249 : AOI21D0BWP7T port map(A1 => n_230, A2 => n_172, B => n_258, ZN => n_231);
  g25227 : ND2D0BWP7T port map(A1 => n_229, A2 => n_327, ZN => n_301);
  g25212 : IND3D0BWP7T port map(A1 => n_264, B1 => n_139, B2 => n_234, ZN => n_372);
  g25242 : NR2XD0BWP7T port map(A1 => n_228, A2 => counter(2), ZN => n_254);
  g25228 : IND2D0BWP7T port map(A1 => n_302, B1 => counter(3), ZN => n_419);
  g25230 : NR2D0BWP7T port map(A1 => n_262, A2 => counter(1), ZN => n_364);
  g25237 : OR2D1BWP7T port map(A1 => n_228, A2 => n_227, Z => n_564);
  g25178 : OR2D1BWP7T port map(A1 => n_574, A2 => n_258, Z => n_645);
  g25176 : ND2D1BWP7T port map(A1 => n_170, A2 => n_268, ZN => n_635);
  g25174 : OR2D1BWP7T port map(A1 => n_574, A2 => n_358, Z => n_549);
  g25172 : OR2D1BWP7T port map(A1 => n_574, A2 => n_255, Z => n_610);
  g25180 : OR2D1BWP7T port map(A1 => n_582, A2 => n_258, Z => n_613);
  g25191 : AOI22D0BWP7T port map(A1 => n_225, A2 => n_93, B1 => n_361, B2 => n_271, ZN => n_226);
  g25130 : INR2XD0BWP7T port map(A1 => n_223, B1 => n_113, ZN => n_224);
  g25132 : NR4D0BWP7T port map(A1 => n_127, A2 => n_72, A3 => n_76, A4 => n_9, ZN => n_222);
  g25146 : AOI22D0BWP7T port map(A1 => n_129, A2 => y(1), B1 => n_488, B2 => sqi_address(1), ZN => n_221);
  g25205 : AOI32D0BWP7T port map(A1 => n_197, A2 => n_242, A3 => counter(1), B1 => n_189, B2 => n_206, ZN => n_219);
  g25204 : AO22D0BWP7T port map(A1 => n_293, A2 => row_buf(0), B1 => edit_buf_in(0), B2 => n_294, Z => n_218);
  g25163 : NR3D0BWP7T port map(A1 => n_171, A2 => y(1), A3 => y(2), ZN => n_217);
  g25165 : AOI21D0BWP7T port map(A1 => n_215, A2 => n_83, B => y(4), ZN => n_216);
  g25186 : AO21D0BWP7T port map(A1 => n_164, A2 => y(2), B => n_213, Z => n_214);
  g25120 : AOI32D0BWP7T port map(A1 => n_459, A2 => n_246, A3 => n_211, B1 => n_150, B2 => y(7), ZN => n_212);
  g25195 : MAOI22D0BWP7T port map(A1 => n_209, A2 => n_118, B1 => n_208, B2 => n_86, ZN => n_210);
  g25196 : OAI211D0BWP7T port map(A1 => n_271, A2 => n_206, B => n_225, C => n_327, ZN => n_207);
  g25199 : MAOI22D0BWP7T port map(A1 => n_124, A2 => n_204, B1 => n_203, B2 => n_245, ZN => n_205);
  g25200 : AOI32D0BWP7T port map(A1 => n_668, A2 => n_410, A3 => n_358, B1 => n_488, B2 => sqi_address(13), ZN => n_202);
  g25202 : AOI32D0BWP7T port map(A1 => n_319, A2 => n_143, A3 => state(0), B1 => n_195, B2 => state(1), ZN => n_200);
  g25203 : AO22D0BWP7T port map(A1 => n_294, A2 => edit_buf_in(7), B1 => calc_buf_in(1), B2 => n_293, Z => n_199);
  g25152 : INVD1BWP7T port map(I => n_343, ZN => n_338);
  g25151 : INVD1BWP7T port map(I => n_345, ZN => n_341);
  g25255 : OA211D0BWP7T port map(A1 => n_504, A2 => n_246, B => n_197, C => n_393, Z => n_198);
  g25209 : AOI22D0BWP7T port map(A1 => n_195, A2 => state(2), B1 => n_152, B2 => n_22, ZN => n_196);
  g25293 : AOI21D0BWP7T port map(A1 => n_192, A2 => counter(0), B => n_230, ZN => n_194);
  g25292 : AOI21D0BWP7T port map(A1 => n_255, A2 => n_192, B => n_142, ZN => n_193);
  g25219 : AOI21D0BWP7T port map(A1 => n_187, A2 => n_132, B => n_197, ZN => n_191);
  g25220 : OAI21D0BWP7T port map(A1 => n_189, A2 => n_180, B => n_105, ZN => n_190);
  g25266 : AOI22D0BWP7T port map(A1 => n_366, A2 => n_185, B1 => n_187, B2 => n_50, ZN => n_188);
  g25244 : IND3D0BWP7T port map(A1 => y(7), B1 => n_185, B2 => n_361, ZN => n_186);
  g25248 : OAI211D0BWP7T port map(A1 => n_242, A2 => n_44, B => n_225, C => n_183, ZN => n_184);
  g25206 : OAI33D0BWP7T port map(A1 => n_178, A2 => n_168, A3 => n_256, B1 => counter(6), B2 => n_227, B3 => n_177, ZN => n_182);
  g25256 : AOI22D0BWP7T port map(A1 => n_180, A2 => n_271, B1 => n_366, B2 => counter(6), ZN => n_181);
  g25259 : MAOI22D0BWP7T port map(A1 => n_189, A2 => n_178, B1 => n_51, B2 => n_177, ZN => n_179);
  g25263 : MAOI22D0BWP7T port map(A1 => n_36, A2 => n_175, B1 => n_203, B2 => n_252, ZN => n_176);
  g25264 : AO22D0BWP7T port map(A1 => n_119, A2 => n_237, B1 => n_178, B2 => n_366, Z => n_174);
  g25265 : MOAI22D0BWP7T port map(A1 => n_172, A2 => n_13, B1 => n_366, B2 => n_242, ZN => n_173);
  g25213 : ND3D0BWP7T port map(A1 => n_171, A2 => n_131, A3 => n_145, ZN => n_277);
  g25217 : INVD1BWP7T port map(I => n_170, ZN => n_597);
  g25239 : ND2D1BWP7T port map(A1 => n_1820, A2 => counter(2), ZN => n_561);
  g25208 : OAI22D0BWP7T port map(A1 => n_100, A2 => n_321, B1 => n_168, B2 => counter(3), ZN => n_169);
  g25224 : IND2D0BWP7T port map(A1 => n_280, B1 => n_183, ZN => n_167);
  g25190 : OA21D0BWP7T port map(A1 => n_134, A2 => n_90, B => n_319, Z => n_166);
  g25187 : AO21D0BWP7T port map(A1 => n_164, A2 => y(4), B => n_163, Z => n_165);
  g25168 : OA21D0BWP7T port map(A1 => n_244, A2 => n_178, B => n_247, Z => n_279);
  g25211 : OA21D0BWP7T port map(A1 => n_244, A2 => n_162, B => n_247, Z => n_238);
  g25135 : OAI221D0BWP7T port map(A1 => n_125, A2 => state(3), B1 => state(2), B2 => n_319, C => n_101, ZN => n_236);
  g25215 : IND3D0BWP7T port map(A1 => n_280, B1 => counter(4), B2 => n_162, ZN => n_380);
  g25183 : NR2XD0BWP7T port map(A1 => n_161, A2 => n_255, ZN => n_343);
  g25182 : NR2XD0BWP7T port map(A1 => n_161, A2 => n_245, ZN => n_345);
  g25169 : NR4D0BWP7T port map(A1 => n_88, A2 => n_30, A3 => n_160, A4 => n_21, ZN => n_239);
  g25232 : OR2D1BWP7T port map(A1 => n_157, A2 => n_321, Z => n_582);
  g25233 : OR2D1BWP7T port map(A1 => n_436, A2 => n_255, Z => n_455);
  g25234 : OR2D1BWP7T port map(A1 => n_436, A2 => n_358, Z => n_470);
  g25246 : ND3D0BWP7T port map(A1 => n_189, A2 => n_369, A3 => n_242, ZN => n_159);
  g25302 : AOI21D0BWP7T port map(A1 => n_141, A2 => counter(3), B => n_375, ZN => n_257);
  g25275 : INR2D0BWP7T port map(A1 => n_158, B1 => counter(4), ZN => n_229);
  g25274 : ND2D0BWP7T port map(A1 => n_158, A2 => n_183, ZN => n_371);
  g25241 : NR2XD0BWP7T port map(A1 => n_157, A2 => n_156, ZN => n_170);
  g25307 : INVD0BWP7T port map(I => n_155, ZN => n_269);
  g25269 : INVD0BWP7T port map(I => n_1820, ZN => n_228);
  g25278 : ND2D0BWP7T port map(A1 => n_209, A2 => counter(6), ZN => n_302);
  g25281 : ND2D0BWP7T port map(A1 => n_209, A2 => n_393, ZN => n_264);
  g25283 : NR2D0BWP7T port map(A1 => n_197, A2 => n_187, ZN => n_262);
  g25236 : OR2D1BWP7T port map(A1 => n_429, A2 => n_258, Z => n_444);
  g25238 : OR2D1BWP7T port map(A1 => n_429, A2 => n_255, Z => n_477);
  g25235 : OR2D1BWP7T port map(A1 => n_429, A2 => n_358, Z => n_473);
  g25240 : OR2D1BWP7T port map(A1 => n_157, A2 => n_309, Z => n_574);
  g25160 : OAI31D0BWP7T port map(A1 => state(0), A2 => n_89, A3 => n_152, B => n_92, ZN => n_153);
  g25184 : INVD0BWP7T port map(I => n_150, ZN => n_151);
  g25247 : MAOI22D0BWP7T port map(A1 => n_74, A2 => n_49, B1 => n_147, B2 => n_255, ZN => n_148);
  g25223 : OAI21D0BWP7T port map(A1 => n_140, A2 => state(0), B => state(1), ZN => n_146);
  g25226 : OAI21D0BWP7T port map(A1 => n_126, A2 => n_145, B => n_103, ZN => n_213);
  g25216 : MOAI22D1BWP7T port map(A1 => n_144, A2 => n_143, B1 => n_84, B2 => state(0), ZN => n_295);
  g25093 : NR4D1BWP7T port map(A1 => n_82, A2 => n_23, A3 => n_46, A4 => n_143, ZN => n_359);
  g25310 : INVD0BWP7T port map(I => n_209, ZN => n_142);
  g25304 : IND3D0BWP7T port map(A1 => y(3), B1 => n_204, B2 => n_85, ZN => n_171);
  g25271 : INVD0BWP7T port map(I => n_386, ZN => n_388);
  g25318 : ND2D0BWP7T port map(A1 => n_141, A2 => n_355, ZN => n_155);
  g25332 : INVD0BWP7T port map(I => n_189, ZN => n_377);
  g25267 : OA22D0BWP7T port map(A1 => n_140, A2 => n_273, B1 => rw, B2 => n_81, Z => n_223);
  g25289 : INVD0BWP7T port map(I => n_500, ZN => n_493);
  g25344 : ND2D0BWP7T port map(A1 => n_141, A2 => n_139, ZN => n_230);
  g25245 : ND3D0BWP7T port map(A1 => n_137, A2 => n_273, A3 => n_136, ZN => n_138);
  g25166 : OAI211D0BWP7T port map(A1 => y(7), A2 => n_134, B => n_130, C => n_211, ZN => n_135);
  g25161 : OAI211D0BWP7T port map(A1 => n_132, A2 => n_134, B => n_131, C => n_130, ZN => n_133);
  g25222 : AO21D0BWP7T port map(A1 => n_164, A2 => y(0), B => n_128, Z => n_129);
  g25257 : OAI22D0BWP7T port map(A1 => n_112, A2 => n_48, B1 => n_152, B2 => n_73, ZN => n_127);
  g25210 : OAI21D0BWP7T port map(A1 => n_126, A2 => n_130, B => n_78, ZN => n_150);
  g25229 : ND2D1BWP7T port map(A1 => n_125, A2 => n_56, ZN => n_161);
  g25268 : INVD0BWP7T port map(I => n_124, ZN => n_215);
  g25276 : INR2D0BWP7T port map(A1 => n_140, B1 => state(0), ZN => n_195);
  g25225 : AO21D0BWP7T port map(A1 => n_164, A2 => n_61, B => n_128, Z => n_163);
  g25277 : ND2D1BWP7T port map(A1 => n_123, A2 => counter(4), ZN => n_157);
  g25231 : AOI211D0BWP7T port map(A1 => n_325, A2 => n_110, B => n_131, C => n_19, ZN => n_247);
  g25284 : IND2D0BWP7T port map(A1 => n_137, B1 => sqi_finished, ZN => n_280);
  g25285 : ND2D1BWP7T port map(A1 => n_123, A2 => n_122, ZN => n_386);
  g25286 : OA21D0BWP7T port map(A1 => n_58, A2 => n_121, B => edit, Z => n_294);
  g25287 : ND2D1BWP7T port map(A1 => n_123, A2 => n_120, ZN => n_436);
  g25340 : OAI21D0BWP7T port map(A1 => n_311, A2 => n_258, B => n_208, ZN => n_119);
  g25296 : OAI22D0BWP7T port map(A1 => n_369, A2 => counter(3), B1 => n_245, B2 => n_321, ZN => n_118);
  g25291 : IND3D0BWP7T port map(A1 => n_147, B1 => counter(1), B2 => n_183, ZN => n_117);
  g25315 : IND2D0BWP7T port map(A1 => n_177, B1 => n_327, ZN => n_172);
  g25314 : NR2D0BWP7T port map(A1 => n_116, A2 => n_47, ZN => n_180);
  g25316 : NR2D0BWP7T port map(A1 => n_208, A2 => counter(6), ZN => n_158);
  g25317 : NR2D0BWP7T port map(A1 => n_116, A2 => counter(7), ZN => n_668);
  g25319 : NR2D0BWP7T port map(A1 => n_116, A2 => counter(2), ZN => n_187);
  g25321 : IND2D0BWP7T port map(A1 => n_147, B1 => y(6), ZN => n_203);
  g25325 : NR2D0BWP7T port map(A1 => n_314, A2 => n_115, ZN => n_197);
  g25323 : NR2D0BWP7T port map(A1 => n_314, A2 => n_504, ZN => n_225);
  g25346 : NR2D0BWP7T port map(A1 => n_314, A2 => n_156, ZN => n_361);
  g25328 : NR2D0BWP7T port map(A1 => n_314, A2 => n_242, ZN => n_209);
  g25350 : NR2D0BWP7T port map(A1 => n_314, A2 => n_309, ZN => n_189);
  g25306 : ND3D0BWP7T port map(A1 => n_114, A2 => n_87, A3 => n_122, ZN => n_500);
  g25288 : ND2D1BWP7T port map(A1 => n_123, A2 => n_237, ZN => n_429);
  g25198 : OAI222D0BWP7T port map(A1 => n_112, A2 => n_111, B1 => n_110, B2 => n_71, C1 => sqi_finished, C2 => n_109, ZN => n_113);
  new_row_buf_reg_5 : LNQD1BWP7T port map(D => n_69, EN => n_108, Q => new_row_buf(5));
  new_row_buf_reg_1 : LNQD1BWP7T port map(D => n_65, EN => n_108, Q => new_row_buf(1));
  new_row_buf_reg_3 : LNQD1BWP7T port map(D => n_68, EN => n_108, Q => new_row_buf(3));
  new_row_buf_reg_0 : LNQD1BWP7T port map(D => n_66, EN => n_108, Q => new_row_buf(0));
  g25192 : IND4D0BWP7T port map(A1 => n_106, B1 => n_204, B2 => n_120, B3 => n_105, ZN => n_107);
  new_row_buf_reg_4 : LNQD1BWP7T port map(D => n_63, EN => n_108, Q => new_row_buf(4));
  g25270 : INVD0BWP7T port map(I => n_128, ZN => n_103);
  g25273 : ND2D0BWP7T port map(A1 => n_152, A2 => n_101, ZN => n_102);
  g25290 : OA21D0BWP7T port map(A1 => n_258, A2 => n_393, B => n_99, Z => n_100);
  g25279 : INR2D0BWP7T port map(A1 => n_134, B1 => n_106, ZN => n_124);
  g25295 : AOI22D0BWP7T port map(A1 => n_175, A2 => n_31, B1 => n_488, B2 => sqi_address(7), ZN => n_97);
  g25297 : AOI22D0BWP7T port map(A1 => n_175, A2 => n_8, B1 => n_488, B2 => sqi_address(6), ZN => n_95);
  g25298 : OAI22D0BWP7T port map(A1 => n_42, A2 => n_168, B1 => n_27, B2 => counter(6), ZN => n_93);
  g25299 : AOI22D0BWP7T port map(A1 => n_307, A2 => n_131, B1 => n_53, B2 => sqi_finished, ZN => n_92);
  g25300 : OAI22D0BWP7T port map(A1 => n_43, A2 => n_358, B1 => n_115, B2 => counter(1), ZN => n_91);
  g25294 : AOI21D0BWP7T port map(A1 => n_204, A2 => n_45, B => n_89, ZN => n_90);
  g25311 : NR2D0BWP7T port map(A1 => n_87, A2 => state(3), ZN => n_88);
  new_row_buf_reg_2 : LNQD1BWP7T port map(D => n_64, EN => n_108, Q => new_row_buf(2));
  g25338 : AOI21D0BWP7T port map(A1 => n_237, A2 => n_258, B => n_62, ZN => n_86);
  g25355 : INVD0BWP7T port map(I => n_314, ZN => n_141);
  g25324 : ND2D0BWP7T port map(A1 => n_409, A2 => counter(2), ZN => n_256);
  g25308 : INVD0BWP7T port map(I => n_134, ZN => n_85);
  g25301 : OAI22D0BWP7T port map(A1 => n_33, A2 => edit, B1 => n_319, B2 => state(1), ZN => n_84);
  g25272 : OR2D0BWP7T port map(A1 => n_106, A2 => n_39, Z => n_83);
  g25162 : OAI211D0BWP7T port map(A1 => n_111, A2 => state(3), B => n_14, C => n_81, ZN => n_82);
  g25303 : NR3D0BWP7T port map(A1 => n_77, A2 => n_55, A3 => state(2), ZN => n_125);
  g25313 : NR2D0BWP7T port map(A1 => n_80, A2 => counter(6), ZN => n_206);
  g25312 : OAI21D0BWP7T port map(A1 => n_268, A2 => n_18, B => n_175, ZN => n_232);
  g25320 : INR2D0BWP7T port map(A1 => n_79, B1 => n_114, ZN => n_137);
  g25282 : ND2D0BWP7T port map(A1 => n_78, A2 => n_311, ZN => n_128);
  g25327 : NR2XD0BWP7T port map(A1 => n_77, A2 => n_79, ZN => n_123);
  g25335 : OAI22D0BWP7T port map(A1 => n_144, A2 => n_110, B1 => n_81, B2 => mode, ZN => n_76);
  g25337 : OAI22D0BWP7T port map(A1 => n_168, A2 => n_227, B1 => n_25, B2 => n_242, ZN => n_75);
  g25334 : OAI21D0BWP7T port map(A1 => n_28, A2 => n_73, B => n_126, ZN => n_74);
  g25333 : AOI21D0BWP7T port map(A1 => n_71, A2 => n_136, B => sqi_finished, ZN => n_72);
  g25363 : ND2D0BWP7T port map(A1 => n_175, A2 => n_70, ZN => n_177);
  g25345 : INR2XD0BWP7T port map(A1 => n_105, B1 => n_307, ZN => n_140);
  g25364 : IND2D0BWP7T port map(A1 => y(7), B1 => n_175, ZN => n_147);
  g25366 : ND2D0BWP7T port map(A1 => n_175, A2 => counter(5), ZN => n_208);
  g25375 : INVD0BWP7T port map(I => n_409, ZN => n_116);
  g25354 : INVD0BWP7T port map(I => n_325, ZN => n_244);
  g25371 : ND2D0BWP7T port map(A1 => n_175, A2 => counter(4), ZN => n_314);
  g25254 : MOAI22D0BWP7T port map(A1 => n_136, A2 => n_648, B1 => n_67, B2 => row_buf(5), ZN => n_69);
  g25243 : MOAI22D0BWP7T port map(A1 => n_136, A2 => n_653, B1 => n_67, B2 => row_buf(3), ZN => n_68);
  g25250 : MOAI22D0BWP7T port map(A1 => n_136, A2 => n_2, B1 => n_67, B2 => row_buf(0), ZN => n_66);
  g25251 : MOAI22D0BWP7T port map(A1 => n_136, A2 => n_1, B1 => n_67, B2 => row_buf(1), ZN => n_65);
  g25252 : MOAI22D0BWP7T port map(A1 => n_136, A2 => n_641, B1 => n_67, B2 => row_buf(2), ZN => n_64);
  g25253 : MOAI22D0BWP7T port map(A1 => n_136, A2 => n_650, B1 => n_67, B2 => row_buf(4), ZN => n_63);
  g25353 : INVD0BWP7T port map(I => n_307, ZN => n_62);
  g25305 : NR3D0BWP7T port map(A1 => n_61, A2 => y(5), A3 => y(4), ZN => n_130);
  g25331 : CKND1BWP7T port map(I => n_60, ZN => n_152);
  g25326 : ND2D1BWP7T port map(A1 => n_122, A2 => n_105, ZN => n_134);
  g25341 : IOA21D0BWP7T port map(A1 => n_227, A2 => counter(6), B => n_324, ZN => n_59);
  g25356 : NR2D0BWP7T port map(A1 => n_144, A2 => state(1), ZN => n_58);
  g25339 : AOI21D0BWP7T port map(A1 => n_418, A2 => n_327, B => n_7, ZN => n_57);
  g25342 : IAO21D0BWP7T port map(A1 => n_234, A2 => counter(6), B => n_271, ZN => n_99);
  g25352 : CKND1BWP7T port map(I => n_77, ZN => n_87);
  g25362 : INR2D0BWP7T port map(A1 => y(7), B1 => n_311, ZN => n_459);
  g25392 : NR2D0BWP7T port map(A1 => n_311, A2 => n_240, ZN => n_409);
  g25370 : IND2D0BWP7T port map(A1 => n_56, B1 => n_79, ZN => n_325);
  g25374 : INVD0BWP7T port map(I => n_80, ZN => n_369);
  g25365 : INR2D0BWP7T port map(A1 => n_237, B1 => n_311, ZN => n_375);
  g25391 : NR2D0BWP7T port map(A1 => n_311, A2 => n_55, ZN => n_366);
  g25357 : IND2D0BWP7T port map(A1 => n_53, B1 => n_136, ZN => n_54);
  g25385 : ND2D5BWP7T port map(A1 => n_17, A2 => n_320, ZN => ready);
  g25336 : AOI32D0BWP7T port map(A1 => n_50, A2 => n_355, A3 => n_49, B1 => n_268, B2 => counter(2), ZN => n_51);
  g25330 : INVD0BWP7T port map(I => n_111, ZN => n_48);
  g25348 : OAI31D0BWP7T port map(A1 => n_70, A2 => n_327, A3 => n_47, B => n_105, ZN => n_60);
  g25343 : AOI221D0BWP7T port map(A1 => n_46, A2 => state(0), B1 => n_16, B2 => state(3), C => n_121, ZN => n_78);
  g25322 : ND2D0BWP7T port map(A1 => n_131, A2 => n_45, ZN => n_106);
  g25329 : NR2D1BWP7T port map(A1 => n_20, A2 => state(2), ZN => n_293);
  g25444 : INVD0BWP7T port map(I => n_311, ZN => n_175);
  g25358 : NR2D0BWP7T port map(A1 => n_418, A2 => n_393, ZN => n_44);
  g25384 : AOI21D0BWP7T port map(A1 => n_139, A2 => n_34, B => n_183, ZN => n_43);
  g25383 : OA21D0BWP7T port map(A1 => n_268, A2 => n_327, B => n_115, Z => n_42);
  g25381 : OAI21D0BWP7T port map(A1 => n_255, A2 => counter(2), B => n_227, ZN => n_41);
  g25360 : NR2D0BWP7T port map(A1 => n_227, A2 => n_327, ZN => n_162);
  g25361 : AN2D1BWP7T port map(A1 => n_56, A2 => n_89, Z => n_114);
  g25367 : ND2D1BWP7T port map(A1 => n_105, A2 => sqi_finished, ZN => n_77);
  g25390 : ND2D0BWP7T port map(A1 => n_40, A2 => n_258, ZN => n_80);
  g25369 : INR2XD0BWP7T port map(A1 => n_39, B1 => y(4), ZN => n_204);
  g25368 : ND2D1BWP7T port map(A1 => n_120, A2 => n_358, ZN => n_307);
  g25382 : OAI22D0BWP7T port map(A1 => n_245, A2 => counter(5), B1 => n_358, B2 => n_242, ZN => n_38);
  g25380 : ND3D0BWP7T port map(A1 => n_131, A2 => n_145, A3 => y(2), ZN => n_37);
  g25379 : OAI21D0BWP7T port map(A1 => n_245, A2 => y(6), B => n_255, ZN => n_36);
  g25377 : MAOI22D0BWP7T port map(A1 => counter(0), A2 => n_34, B1 => n_245, B2 => n_49, ZN => n_35);
  g25376 : AOI21D0BWP7T port map(A1 => n_160, A2 => n_319, B => n_46, ZN => n_33);
  g25378 : OAI22D0BWP7T port map(A1 => n_309, A2 => n_246, B1 => n_115, B2 => counter(0), ZN => n_32);
  g25359 : OAI21D0BWP7T port map(A1 => n_4, A2 => n_46, B => state(0), ZN => n_112);
  g25393 : INVD0BWP7T port map(I => n_31, ZN => n_192);
  g25387 : AOI22D0BWP7T port map(A1 => n_30, A2 => n_24, B1 => n_46, B2 => FE_OFN2_n_0, ZN => n_286);
  g25373 : INVD0BWP7T port map(I => n_45, ZN => n_61);
  g25347 : AOI21D0BWP7T port map(A1 => n_5, A2 => n_3, B => edit, ZN => n_111);
  g25389 : NR2XD0BWP7T port map(A1 => n_55, A2 => n_258, ZN => n_122);
  g25351 : NR3D0BWP7T port map(A1 => n_136, A2 => state(2), A3 => sqi_finished, ZN => n_108);
  g25473 : ND2D1BWP7T port map(A1 => n_50, A2 => sqi_data_in(2), ZN => n_596);
  g25372 : ND2D0BWP7T port map(A1 => n_136, A2 => n_29, ZN => n_488);
  g25448 : NR2D0BWP7T port map(A1 => n_268, A2 => n_178, ZN => n_28);
  g25447 : NR2D0BWP7T port map(A1 => n_183, A2 => n_139, ZN => n_27);
  g25442 : INVD0BWP7T port map(I => n_418, ZN => n_26);
  g25450 : NR2D0BWP7T port map(A1 => n_268, A2 => n_393, ZN => n_25);
  g25430 : NR2D0BWP7T port map(A1 => n_24, A2 => n_81, ZN => n_250);
  g25433 : ND2D1BWP7T port map(A1 => n_23, A2 => state(1), ZN => n_71);
  g25456 : ND2D1BWP7T port map(A1 => n_22, A2 => n_319, ZN => n_109);
  g25457 : NR2D0BWP7T port map(A1 => n_268, A2 => n_355, ZN => n_363);
  g25439 : ND2D1BWP7T port map(A1 => n_23, A2 => state(0), ZN => n_144);
  g25458 : ND2D1BWP7T port map(A1 => n_22, A2 => state(0), ZN => n_79);
  g25461 : ND2D1BWP7T port map(A1 => n_50, A2 => sqi_data_in(6), ZN => n_625);
  g25462 : ND2D1BWP7T port map(A1 => n_50, A2 => sqi_data_in(7), ZN => n_578);
  g25470 : ND2D1BWP7T port map(A1 => n_50, A2 => sqi_data_in(3), ZN => n_592);
  g25466 : ND2D1BWP7T port map(A1 => n_50, A2 => sqi_data_in(4), ZN => n_590);
  g25471 : ND2D1BWP7T port map(A1 => n_50, A2 => sqi_data_in(5), ZN => n_587);
  g25476 : ND2D1BWP7T port map(A1 => n_22, A2 => n_21, ZN => n_311);
  g25386 : AOI22D0BWP7T port map(A1 => n_21, A2 => state(1), B1 => n_101, B2 => state(3), ZN => n_20);
  g25394 : INVD0BWP7T port map(I => n_73, ZN => n_19);
  g25395 : INR2D0BWP7T port map(A1 => n_49, B1 => counter(1), ZN => n_18);
  g25451 : ND2D1BWP7T port map(A1 => n_30, A2 => state(1), ZN => n_17);
  g25437 : NR2D0BWP7T port map(A1 => n_246, A2 => n_132, ZN => n_31);
  g25410 : INVD5BWP7T port map(I => n_692, ZN => sqi_address(10));
  g25429 : INVD5BWP7T port map(I => n_685, ZN => sqi_address(11));
  g25408 : INVD5BWP7T port map(I => n_693, ZN => sqi_address(9));
  g25404 : INVD5BWP7T port map(I => n_695, ZN => sqi_address(12));
  g25398 : INVD5BWP7T port map(I => n_698, ZN => sqi_address(7));
  g25400 : INVD5BWP7T port map(I => n_697, ZN => sqi_address(4));
  g25402 : INVD5BWP7T port map(I => n_696, ZN => sqi_address(6));
  g25406 : INVD5BWP7T port map(I => n_694, ZN => sqi_address(3));
  g25388 : INR3D0BWP7T port map(A1 => n_145, B1 => y(3), B2 => y(2), ZN => n_45);
  g25443 : INVD1BWP7T port map(I => n_131, ZN => n_273);
  g25441 : CKND1BWP7T port map(I => n_55, ZN => n_120);
  g25349 : IND4D0BWP7T port map(A1 => n_16, B1 => n_15, B2 => state(3), B3 => n_126, ZN => n_67);
  g25467 : ND2D1BWP7T port map(A1 => n_255, A2 => n_319, ZN => n_401);
  g25415 : INVD5BWP7T port map(I => n_690, ZN => sqi_address(14));
  g25417 : INVD5BWP7T port map(I => n_689, ZN => sqi_address(8));
  g25419 : INVD5BWP7T port map(I => n_688, ZN => sqi_address(2));
  g25421 : INVD5BWP7T port map(I => n_687, ZN => sqi_address(1));
  g25427 : INVD5BWP7T port map(I => n_686, ZN => sqi_address(0));
  g25432 : INVD5BWP7T port map(I => n_684, ZN => sqi_address(13));
  g25434 : NR2XD0BWP7T port map(A1 => n_132, A2 => y(5), ZN => n_39);
  g25436 : NR2D0BWP7T port map(A1 => n_29, A2 => n_101, ZN => n_53);
  g25453 : IND2D0BWP7T port map(A1 => n_49, B1 => n_246, ZN => n_40);
  g25413 : INVD5BWP7T port map(I => n_691, ZN => sqi_address(5));
  g25455 : NR2XD0BWP7T port map(A1 => n_14, A2 => state(1), ZN => n_56);
  g25459 : ND2D0BWP7T port map(A1 => n_178, A2 => n_132, ZN => n_234);
  g25464 : NR2XD0BWP7T port map(A1 => n_156, A2 => counter(4), ZN => n_237);
  g25463 : ND2D1BWP7T port map(A1 => n_258, A2 => n_319, ZN => n_403);
  g25465 : NR2XD0BWP7T port map(A1 => n_13, A2 => counter(7), ZN => n_105);
  g25469 : AOI21D0BWP7T port map(A1 => counter(1), A2 => y(7), B => n_178, ZN => n_418);
  g25472 : ND2D1BWP7T port map(A1 => n_178, A2 => counter(2), ZN => n_227);
  g25474 : ND2D1BWP7T port map(A1 => n_245, A2 => n_319, ZN => n_405);
  sqi_address_reg_9 : DFKCND1BWP7T port map(CN => new_sqi_address(9), CP => CTS_14, D => FE_OFN2_n_0, Q => UNCONNECTED9, QN => n_693);
  g25449 : AOI21D0BWP7T port map(A1 => n_143, A2 => sqi_finished, B => state(2), ZN => n_12);
  sqi_address_reg_5 : DFKCND1BWP7T port map(CN => new_sqi_address(5), CP => CTS_14, D => FE_OFN1_n_0, Q => UNCONNECTED10, QN => n_691);
  sqi_address_reg_4 : DFKCND1BWP7T port map(CN => new_sqi_address(4), CP => CTS_14, D => FE_OFN1_n_0, Q => UNCONNECTED11, QN => n_697);
  sqi_address_reg_8 : DFKCND1BWP7T port map(CN => new_sqi_address(8), CP => CTS_14, D => FE_OFN2_n_0, Q => UNCONNECTED12, QN => n_689);
  sqi_address_reg_12 : DFKCND1BWP7T port map(CN => new_sqi_address(12), CP => CTS_14, D => FE_OFN3_n_0, Q => UNCONNECTED13, QN => n_695);
  sqi_address_reg_7 : DFKCND1BWP7T port map(CN => new_sqi_address(7), CP => CTS_14, D => FE_OFN1_n_0, Q => UNCONNECTED14, QN => n_698);
  sqi_address_reg_1 : DFKCND1BWP7T port map(CN => new_sqi_address(1), CP => CTS_14, D => FE_OFN1_n_0, Q => UNCONNECTED15, QN => n_687);
  sqi_address_reg_0 : DFKCND1BWP7T port map(CN => new_sqi_address(0), CP => CTS_14, D => FE_OFN1_n_0, Q => UNCONNECTED16, QN => n_686);
  sqi_address_reg_6 : DFKCND1BWP7T port map(CN => new_sqi_address(6), CP => CTS_14, D => FE_OFN1_n_0, Q => UNCONNECTED17, QN => n_696);
  sqi_address_reg_14 : DFKCND1BWP7T port map(CN => new_sqi_address(14), CP => CTS_14, D => FE_OFN3_n_0, Q => UNCONNECTED18, QN => n_690);
  g25396 : NR2D0BWP7T port map(A1 => n_10, A2 => ce, ZN => n_11);
  g25505 : INVD0BWP7T port map(I => n_255, ZN => n_185);
  row_buf_reg_2 : DFKCNQD1BWP7T port map(CN => new_row_buf(2), CP => CTS_13, D => FE_OFN2_n_0, Q => row_buf(2));
  row_buf_reg_4 : DFKCNQD1BWP7T port map(CN => new_row_buf(4), CP => CTS_13, D => n_0, Q => row_buf(4));
  row_buf_reg_0 : DFKCNQD1BWP7T port map(CN => new_row_buf(0), CP => CTS_13, D => FE_OFN2_n_0, Q => row_buf(0));
  g25438 : ND2D1BWP7T port map(A1 => n_21, A2 => state(2), ZN => n_73);
  g25501 : INVD0BWP7T port map(I => n_321, ZN => n_139);
  g25479 : INVD0BWP7T port map(I => n_13, ZN => n_271);
  g25460 : CKND2D1BWP7T port map(A1 => n_319, A2 => n_358, ZN => n_400);
  g25507 : INVD1BWP7T port map(I => n_258, ZN => n_268);
  sqi_address_reg_10 : DFKCND1BWP7T port map(CN => new_sqi_address(10), CP => CTS_14, D => FE_OFN3_n_0, Q => UNCONNECTED19, QN => n_692);
  sqi_address_reg_2 : DFKCND1BWP7T port map(CN => new_sqi_address(2), CP => CTS_14, D => FE_OFN1_n_0, Q => UNCONNECTED20, QN => n_688);
  sqi_address_reg_3 : DFKCND1BWP7T port map(CN => new_sqi_address(3), CP => CTS_14, D => FE_OFN1_n_0, Q => UNCONNECTED21, QN => n_694);
  sqi_address_reg_13 : DFKCND1BWP7T port map(CN => new_sqi_address(13), CP => CTS_14, D => FE_OFN3_n_0, Q => UNCONNECTED22, QN => n_684);
  sqi_address_reg_11 : DFKCND1BWP7T port map(CN => new_sqi_address(11), CP => CTS_14, D => FE_OFN3_n_0, Q => UNCONNECTED23, QN => n_685);
  g25445 : OA21D0BWP7T port map(A1 => state(3), A2 => sqi_finished, B => n_16, Z => n_9);
  g25452 : OAI22D0BWP7T port map(A1 => n_252, A2 => y(6), B1 => counter(0), B2 => n_211, ZN => n_8);
  row_buf_reg_3 : DFKCNQD1BWP7T port map(CN => new_row_buf(3), CP => CTS_13, D => n_0, Q => row_buf(3));
  row_buf_reg_5 : DFKCNQD1BWP7T port map(CN => new_row_buf(5), CP => CTS_13, D => n_0, Q => row_buf(5));
  row_buf_reg_1 : DFKCNQD1BWP7T port map(CN => new_row_buf(1), CP => CTS_13, D => FE_OFN2_n_0, Q => row_buf(1));
  g25454 : NR2D1BWP7T port map(A1 => n_126, A2 => n_15, ZN => n_121);
  g25498 : INVD1BWP7T port map(I => n_29, ZN => n_23);
  g25468 : ND2D1BWP7T port map(A1 => n_7, A2 => n_70, ZN => n_55);
  g25500 : INVD1BWP7T port map(I => n_30, ZN => n_81);
  g25499 : CKND1BWP7T port map(I => n_160, ZN => n_22);
  g25477 : INVD0BWP7T port map(I => n_6, ZN => n_324);
  g25502 : INVD0BWP7T port map(I => n_168, ZN => n_410);
  g25504 : INVD0BWP7T port map(I => n_156, ZN => n_183);
  g25475 : NR2XD0BWP7T port map(A1 => n_126, A2 => state(0), ZN => n_131);
  g25506 : CKND1BWP7T port map(I => n_245, ZN => n_50);
  g25440 : OR2D1BWP7T port map(A1 => n_10, A2 => state(0), Z => n_136);
  g25446 : NR3D0BWP7T port map(A1 => x(3), A2 => x(4), A3 => x(0), ZN => n_5);
  g25508 : NR2D0BWP7T port map(A1 => n_143, A2 => state(3), ZN => n_4);
  g25481 : INVD0BWP7T port map(I => n_126, ZN => n_164);
  g25513 : ND2D1BWP7T port map(A1 => n_143, A2 => state(2), ZN => n_160);
  g25489 : INR2D0BWP7T port map(A1 => y(7), B1 => n_211, ZN => n_49);
  g25516 : ND2D0BWP7T port map(A1 => n_242, A2 => counter(6), ZN => n_168);
  g25478 : INVD1BWP7T port map(I => n_34, ZN => n_132);
  g25482 : CKND1BWP7T port map(I => n_358, ZN => n_178);
  g25480 : INVD1BWP7T port map(I => n_7, ZN => n_309);
  g25520 : ND2D1BWP7T port map(A1 => n_246, A2 => counter(0), ZN => n_245);
  g25497 : INVD0BWP7T port map(I => n_21, ZN => n_14);
  g25491 : NR2D0BWP7T port map(A1 => n_393, A2 => n_242, ZN => n_6);
  g25493 : ND2D1BWP7T port map(A1 => n_242, A2 => n_393, ZN => n_13);
  g25514 : NR2D1BWP7T port map(A1 => n_319, A2 => n_15, ZN => n_30);
  g25510 : ND2D1BWP7T port map(A1 => n_70, A2 => counter(3), ZN => n_240);
  g25512 : ND2D1BWP7T port map(A1 => n_319, A2 => n_89, ZN => n_29);
  g25518 : ND2D1BWP7T port map(A1 => n_327, A2 => counter(2), ZN => n_156);
  g25503 : INVD1BWP7T port map(I => n_320, ZN => n_46);
  g25515 : ND2D1BWP7T port map(A1 => n_355, A2 => counter(3), ZN => n_321);
  g25521 : ND2D1BWP7T port map(A1 => n_252, A2 => n_246, ZN => n_258);
  g25519 : ND2D1BWP7T port map(A1 => n_252, A2 => counter(1), ZN => n_255);
  g25492 : NR2XD0BWP7T port map(A1 => y(6), A2 => y(7), ZN => n_34);
  g25486 : NR2D0BWP7T port map(A1 => state(1), A2 => state(2), ZN => n_16);
  g25494 : NR2XD0BWP7T port map(A1 => counter(2), A2 => counter(3), ZN => n_7);
  g25509 : CKND2D1BWP7T port map(A1 => state(3), A2 => state(1), ZN => n_10);
  g25490 : ND2D0BWP7T port map(A1 => counter(2), A2 => counter(3), ZN => n_115);
  g25511 : NR2D1BWP7T port map(A1 => state(3), A2 => state(0), ZN => n_21);
  g25517 : ND2D1BWP7T port map(A1 => state(3), A2 => state(2), ZN => n_320);
  g25483 : NR2D0BWP7T port map(A1 => x(1), A2 => x(2), ZN => n_3);
  g25484 : NR2D0BWP7T port map(A1 => counter(1), A2 => counter(2), ZN => n_47);
  g25485 : ND2D0BWP7T port map(A1 => state(1), A2 => ce, ZN => n_24);
  g25487 : NR2XD0BWP7T port map(A1 => state(1), A2 => state(0), ZN => n_101);
  g25488 : NR2XD0BWP7T port map(A1 => y(0), A2 => y(1), ZN => n_145);
  g25495 : CKND2D1BWP7T port map(A1 => state(1), A2 => state(2), ZN => n_126);
  g25496 : CKND2D1BWP7T port map(A1 => counter(0), A2 => counter(1), ZN => n_358);
  g25522 : INVD0BWP7T port map(I => sqi_data_in(0), ZN => n_2);
  g25534 : INVD0BWP7T port map(I => y(6), ZN => n_211);
  g25527 : INVD1BWP7T port map(I => sqi_data_in(7), ZN => n_631);
  g25542 : INVD1BWP7T port map(I => sqi_data_in(6), ZN => n_637);
  g25529 : INVD1BWP7T port map(I => sqi_data_in(4), ZN => n_650);
  g25533 : INVD0BWP7T port map(I => sqi_data_in(1), ZN => n_1);
  g25535 : INVD0BWP7T port map(I => sqi_finished, ZN => n_110);
  g25543 : INVD1BWP7T port map(I => sqi_data_in(2), ZN => n_641);
  g25544 : INVD1BWP7T port map(I => sqi_data_in(5), ZN => n_648);
  g25528 : INVD1BWP7T port map(I => sqi_data_in(3), ZN => n_653);
  g25531 : CKND2BWP7T port map(I => reset, ZN => n_0);
  g2 : MAOI22D0BWP7T port map(A1 => n_114, A2 => sqi_finished, B1 => n_60, B2 => n_109, ZN => n_739);
  drc_bufs25799 : INVD5BWP7T port map(I => n_742, ZN => calc_buf_out(2));
  drc_bufs25805 : INVD5BWP7T port map(I => n_748, ZN => framebuffer_buf(157));
  drc_bufs25811 : INVD5BWP7T port map(I => n_754, ZN => framebuffer_buf(156));
  drc_bufs25817 : INVD5BWP7T port map(I => n_760, ZN => framebuffer_buf(155));
  drc_bufs25823 : INVD5BWP7T port map(I => n_766, ZN => framebuffer_buf(154));
  drc_bufs25829 : INVD5BWP7T port map(I => n_772, ZN => framebuffer_buf(153));
  drc_bufs25835 : INVD5BWP7T port map(I => n_778, ZN => framebuffer_buf(152));
  drc_bufs25841 : INVD5BWP7T port map(I => n_784, ZN => framebuffer_buf(151));
  drc_bufs25847 : INVD5BWP7T port map(I => n_790, ZN => framebuffer_buf(150));
  drc_bufs25853 : INVD5BWP7T port map(I => n_796, ZN => framebuffer_buf(149));
  drc_bufs25859 : INVD5BWP7T port map(I => n_802, ZN => framebuffer_buf(148));
  drc_bufs25865 : INVD5BWP7T port map(I => n_808, ZN => framebuffer_buf(147));
  drc_bufs25871 : INVD5BWP7T port map(I => n_814, ZN => framebuffer_buf(146));
  drc_bufs25877 : INVD5BWP7T port map(I => n_820, ZN => framebuffer_buf(145));
  drc_bufs25883 : INVD5BWP7T port map(I => n_826, ZN => framebuffer_buf(144));
  drc_bufs25889 : INVD5BWP7T port map(I => n_832, ZN => framebuffer_buf(143));
  drc_bufs25895 : INVD5BWP7T port map(I => n_838, ZN => framebuffer_buf(142));
  drc_bufs25901 : INVD5BWP7T port map(I => n_844, ZN => framebuffer_buf(141));
  drc_bufs25907 : INVD5BWP7T port map(I => n_850, ZN => framebuffer_buf(140));
  drc_bufs25913 : INVD5BWP7T port map(I => n_856, ZN => framebuffer_buf(139));
  drc_bufs25919 : INVD5BWP7T port map(I => n_862, ZN => framebuffer_buf(138));
  drc_bufs25925 : INVD5BWP7T port map(I => n_868, ZN => calc_buf_out(3));
  drc_bufs25931 : INVD5BWP7T port map(I => n_874, ZN => framebuffer_buf(136));
  drc_bufs25937 : INVD5BWP7T port map(I => n_880, ZN => framebuffer_buf(135));
  drc_bufs25943 : INVD5BWP7T port map(I => n_886, ZN => framebuffer_buf(134));
  drc_bufs25949 : INVD5BWP7T port map(I => n_892, ZN => framebuffer_buf(133));
  drc_bufs25955 : INVD5BWP7T port map(I => n_898, ZN => framebuffer_buf(132));
  drc_bufs25961 : INVD5BWP7T port map(I => n_904, ZN => framebuffer_buf(131));
  drc_bufs25967 : INVD5BWP7T port map(I => n_910, ZN => framebuffer_buf(130));
  drc_bufs25973 : INVD5BWP7T port map(I => n_916, ZN => calc_buf_out(7));
  drc_bufs25979 : INVD5BWP7T port map(I => n_922, ZN => framebuffer_buf(128));
  drc_bufs25985 : INVD5BWP7T port map(I => n_928, ZN => framebuffer_buf(127));
  drc_bufs25991 : INVD5BWP7T port map(I => n_934, ZN => framebuffer_buf(126));
  drc_bufs25997 : INVD5BWP7T port map(I => n_940, ZN => framebuffer_buf(125));
  drc_bufs26003 : INVD5BWP7T port map(I => n_946, ZN => framebuffer_buf(124));
  drc_bufs26009 : INVD5BWP7T port map(I => n_952, ZN => framebuffer_buf(123));
  drc_bufs26015 : INVD5BWP7T port map(I => n_958, ZN => framebuffer_buf(122));
  drc_bufs26021 : INVD5BWP7T port map(I => n_964, ZN => calc_buf_out(15));
  drc_bufs26027 : INVD5BWP7T port map(I => n_970, ZN => framebuffer_buf(120));
  drc_bufs26033 : INVD5BWP7T port map(I => n_976, ZN => framebuffer_buf(119));
  drc_bufs26039 : INVD5BWP7T port map(I => n_982, ZN => framebuffer_buf(118));
  drc_bufs26045 : INVD5BWP7T port map(I => n_988, ZN => framebuffer_buf(115));
  drc_bufs26051 : INVD5BWP7T port map(I => n_994, ZN => framebuffer_buf(114));
  drc_bufs26057 : INVD5BWP7T port map(I => n_1000, ZN => framebuffer_buf(113));
  drc_bufs26063 : INVD5BWP7T port map(I => n_1006, ZN => framebuffer_buf(112));
  drc_bufs26069 : INVD5BWP7T port map(I => n_1012, ZN => framebuffer_buf(7));
  drc_bufs26075 : INVD5BWP7T port map(I => n_1018, ZN => framebuffer_buf(110));
  drc_bufs26081 : INVD5BWP7T port map(I => n_1024, ZN => framebuffer_buf(109));
  drc_bufs26087 : INVD5BWP7T port map(I => n_1030, ZN => framebuffer_buf(108));
  drc_bufs26093 : INVD5BWP7T port map(I => n_1036, ZN => framebuffer_buf(107));
  drc_bufs26099 : INVD5BWP7T port map(I => n_1042, ZN => framebuffer_buf(39));
  drc_bufs26105 : INVD5BWP7T port map(I => n_1048, ZN => framebuffer_buf(103));
  drc_bufs26111 : INVD5BWP7T port map(I => n_1054, ZN => framebuffer_buf(104));
  drc_bufs26117 : INVD5BWP7T port map(I => n_1060, ZN => framebuffer_buf(40));
  drc_bufs26123 : INVD5BWP7T port map(I => n_1066, ZN => framebuffer_buf(102));
  drc_bufs26129 : INVD5BWP7T port map(I => n_1072, ZN => framebuffer_buf(101));
  drc_bufs26135 : INVD5BWP7T port map(I => n_1078, ZN => framebuffer_buf(100));
  drc_bufs26141 : INVD5BWP7T port map(I => n_1084, ZN => framebuffer_buf(99));
  drc_bufs26147 : INVD5BWP7T port map(I => n_1090, ZN => framebuffer_buf(98));
  drc_bufs26153 : INVD5BWP7T port map(I => n_1096, ZN => framebuffer_buf(97));
  drc_bufs26159 : INVD5BWP7T port map(I => n_1102, ZN => framebuffer_buf(96));
  drc_bufs26165 : INVD5BWP7T port map(I => n_1108, ZN => framebuffer_buf(95));
  drc_bufs26171 : INVD5BWP7T port map(I => n_1114, ZN => framebuffer_buf(94));
  drc_bufs26177 : INVD5BWP7T port map(I => n_1120, ZN => framebuffer_buf(93));
  drc_bufs26183 : INVD5BWP7T port map(I => n_1126, ZN => framebuffer_buf(92));
  drc_bufs26189 : INVD5BWP7T port map(I => n_1132, ZN => framebuffer_buf(91));
  drc_bufs26195 : INVD5BWP7T port map(I => n_1138, ZN => framebuffer_buf(90));
  drc_bufs26201 : INVD5BWP7T port map(I => n_1144, ZN => framebuffer_buf(89));
  drc_bufs26207 : INVD5BWP7T port map(I => n_1150, ZN => framebuffer_buf(88));
  drc_bufs26213 : INVD5BWP7T port map(I => n_1156, ZN => framebuffer_buf(87));
  drc_bufs26219 : INVD5BWP7T port map(I => n_1162, ZN => framebuffer_buf(86));
  drc_bufs26225 : INVD5BWP7T port map(I => n_1168, ZN => framebuffer_buf(85));
  drc_bufs26231 : INVD5BWP7T port map(I => n_1174, ZN => framebuffer_buf(84));
  drc_bufs26237 : INVD5BWP7T port map(I => n_1180, ZN => framebuffer_buf(83));
  drc_bufs26243 : INVD5BWP7T port map(I => n_1186, ZN => framebuffer_buf(82));
  drc_bufs26249 : INVD5BWP7T port map(I => n_1192, ZN => framebuffer_buf(81));
  drc_bufs26255 : INVD5BWP7T port map(I => n_1198, ZN => framebuffer_buf(80));
  drc_bufs26261 : INVD5BWP7T port map(I => n_1204, ZN => framebuffer_buf(105));
  drc_bufs26267 : INVD5BWP7T port map(I => n_1210, ZN => framebuffer_buf(78));
  drc_bufs26273 : INVD5BWP7T port map(I => n_1216, ZN => framebuffer_buf(77));
  drc_bufs26279 : INVD5BWP7T port map(I => n_1222, ZN => framebuffer_buf(76));
  drc_bufs26285 : INVD5BWP7T port map(I => n_1228, ZN => framebuffer_buf(106));
  drc_bufs26291 : INVD5BWP7T port map(I => n_1234, ZN => framebuffer_buf(74));
  drc_bufs26297 : INVD5BWP7T port map(I => n_1240, ZN => framebuffer_buf(73));
  drc_bufs26303 : INVD5BWP7T port map(I => n_1246, ZN => framebuffer_buf(72));
  drc_bufs26309 : INVD5BWP7T port map(I => n_1252, ZN => framebuffer_buf(8));
  drc_bufs26315 : INVD5BWP7T port map(I => n_1258, ZN => framebuffer_buf(70));
  drc_bufs26321 : INVD5BWP7T port map(I => n_1264, ZN => framebuffer_buf(69));
  drc_bufs26327 : INVD5BWP7T port map(I => n_1270, ZN => framebuffer_buf(68));
  drc_bufs26333 : INVD5BWP7T port map(I => n_1276, ZN => framebuffer_buf(67));
  drc_bufs26339 : INVD5BWP7T port map(I => n_1282, ZN => framebuffer_buf(66));
  drc_bufs26345 : INVD5BWP7T port map(I => n_1288, ZN => framebuffer_buf(65));
  drc_bufs26351 : INVD5BWP7T port map(I => n_1294, ZN => framebuffer_buf(64));
  drc_bufs26357 : INVD5BWP7T port map(I => n_1300, ZN => framebuffer_buf(63));
  drc_bufs26363 : INVD5BWP7T port map(I => n_1306, ZN => framebuffer_buf(62));
  drc_bufs26369 : INVD5BWP7T port map(I => n_1312, ZN => framebuffer_buf(61));
  drc_bufs26375 : INVD5BWP7T port map(I => n_1318, ZN => framebuffer_buf(60));
  drc_bufs26381 : INVD5BWP7T port map(I => n_1324, ZN => framebuffer_buf(59));
  drc_bufs26387 : INVD5BWP7T port map(I => n_1330, ZN => framebuffer_buf(58));
  drc_bufs26393 : INVD5BWP7T port map(I => n_1336, ZN => framebuffer_buf(57));
  drc_bufs26399 : INVD5BWP7T port map(I => n_1342, ZN => framebuffer_buf(56));
  drc_bufs26405 : INVD5BWP7T port map(I => n_1348, ZN => framebuffer_buf(137));
  drc_bufs26411 : INVD5BWP7T port map(I => n_1354, ZN => framebuffer_buf(54));
  drc_bufs26417 : INVD5BWP7T port map(I => n_1360, ZN => framebuffer_buf(53));
  drc_bufs26423 : INVD5BWP7T port map(I => n_1366, ZN => framebuffer_buf(52));
  drc_bufs26429 : INVD5BWP7T port map(I => n_1372, ZN => framebuffer_buf(129));
  drc_bufs26435 : INVD5BWP7T port map(I => n_1378, ZN => framebuffer_buf(50));
  drc_bufs26441 : INVD5BWP7T port map(I => n_1384, ZN => framebuffer_buf(49));
  drc_bufs26447 : INVD5BWP7T port map(I => n_1390, ZN => framebuffer_buf(48));
  drc_bufs26453 : INVD5BWP7T port map(I => n_1396, ZN => framebuffer_buf(121));
  drc_bufs26459 : INVD5BWP7T port map(I => n_1402, ZN => framebuffer_buf(46));
  drc_bufs26465 : INVD5BWP7T port map(I => n_1408, ZN => framebuffer_buf(45));
  drc_bufs26471 : INVD5BWP7T port map(I => n_1414, ZN => framebuffer_buf(44));
  drc_bufs26477 : INVD5BWP7T port map(I => n_1420, ZN => framebuffer_buf(41));
  drc_bufs26483 : INVD5BWP7T port map(I => n_1426, ZN => framebuffer_buf(42));
  drc_bufs26489 : INVD5BWP7T port map(I => n_1432, ZN => framebuffer_buf(9));
  drc_bufs26495 : INVD5BWP7T port map(I => n_1438, ZN => framebuffer_buf(43));
  drc_bufs26501 : INVD5BWP7T port map(I => n_1444, ZN => framebuffer_buf(111));
  drc_bufs26507 : INVD5BWP7T port map(I => n_1450, ZN => framebuffer_buf(38));
  drc_bufs26513 : INVD5BWP7T port map(I => n_1456, ZN => framebuffer_buf(37));
  drc_bufs26519 : INVD5BWP7T port map(I => n_1462, ZN => framebuffer_buf(36));
  drc_bufs26525 : INVD5BWP7T port map(I => n_1468, ZN => framebuffer_buf(35));
  drc_bufs26531 : INVD5BWP7T port map(I => n_1474, ZN => framebuffer_buf(34));
  drc_bufs26537 : INVD5BWP7T port map(I => n_1480, ZN => framebuffer_buf(33));
  drc_bufs26543 : INVD5BWP7T port map(I => n_1486, ZN => framebuffer_buf(32));
  drc_bufs26549 : INVD5BWP7T port map(I => n_1492, ZN => framebuffer_buf(31));
  drc_bufs26555 : INVD5BWP7T port map(I => n_1498, ZN => framebuffer_buf(30));
  drc_bufs26561 : INVD5BWP7T port map(I => n_1504, ZN => framebuffer_buf(29));
  drc_bufs26567 : INVD5BWP7T port map(I => n_1510, ZN => framebuffer_buf(28));
  drc_bufs26573 : INVD5BWP7T port map(I => n_1516, ZN => framebuffer_buf(79));
  drc_bufs26579 : INVD5BWP7T port map(I => n_1522, ZN => framebuffer_buf(26));
  drc_bufs26585 : INVD5BWP7T port map(I => n_1528, ZN => framebuffer_buf(75));
  drc_bufs26591 : INVD5BWP7T port map(I => n_1534, ZN => framebuffer_buf(24));
  drc_bufs26597 : INVD5BWP7T port map(I => n_1540, ZN => framebuffer_buf(71));
  drc_bufs26603 : INVD5BWP7T port map(I => n_1546, ZN => framebuffer_buf(22));
  drc_bufs26609 : INVD5BWP7T port map(I => n_1552, ZN => framebuffer_buf(21));
  drc_bufs26615 : INVD5BWP7T port map(I => n_1558, ZN => framebuffer_buf(20));
  drc_bufs26621 : INVD5BWP7T port map(I => n_1564, ZN => framebuffer_buf(19));
  drc_bufs26627 : INVD5BWP7T port map(I => n_1570, ZN => framebuffer_buf(18));
  drc_bufs26633 : INVD5BWP7T port map(I => n_1576, ZN => framebuffer_buf(17));
  drc_bufs26639 : INVD5BWP7T port map(I => n_1582, ZN => framebuffer_buf(16));
  drc_bufs26645 : INVD5BWP7T port map(I => n_1588, ZN => framebuffer_buf(55));
  drc_bufs26651 : INVD5BWP7T port map(I => n_1594, ZN => framebuffer_buf(14));
  drc_bufs26657 : INVD5BWP7T port map(I => n_1600, ZN => framebuffer_buf(51));
  drc_bufs26663 : INVD5BWP7T port map(I => n_1606, ZN => framebuffer_buf(12));
  drc_bufs26669 : INVD5BWP7T port map(I => n_1612, ZN => framebuffer_buf(10));
  drc_bufs26675 : INVD5BWP7T port map(I => n_1618, ZN => calc_buf_out(18));
  drc_bufs26681 : INVD5BWP7T port map(I => n_1624, ZN => framebuffer_buf(11));
  drc_bufs26687 : INVD5BWP7T port map(I => n_1630, ZN => framebuffer_buf(47));
  drc_bufs26693 : INVD5BWP7T port map(I => n_1636, ZN => framebuffer_buf(13));
  drc_bufs26699 : INVD5BWP7T port map(I => n_1642, ZN => framebuffer_buf(6));
  drc_bufs26705 : INVD5BWP7T port map(I => n_1648, ZN => framebuffer_buf(5));
  drc_bufs26711 : INVD5BWP7T port map(I => n_1654, ZN => framebuffer_buf(4));
  drc_bufs26717 : INVD5BWP7T port map(I => n_1660, ZN => framebuffer_buf(3));
  drc_bufs26723 : INVD5BWP7T port map(I => n_1666, ZN => framebuffer_buf(2));
  drc_bufs26729 : INVD5BWP7T port map(I => n_1672, ZN => framebuffer_buf(27));
  drc_bufs26735 : INVD5BWP7T port map(I => n_1678, ZN => framebuffer_buf(25));
  drc_bufs26741 : INVD5BWP7T port map(I => n_1684, ZN => framebuffer_buf(23));
  drc_bufs26747 : INVD5BWP7T port map(I => n_1690, ZN => calc_buf_out(22));
  drc_bufs26753 : INVD5BWP7T port map(I => n_1696, ZN => calc_buf_out(21));
  drc_bufs26759 : INVD5BWP7T port map(I => n_1702, ZN => calc_buf_out(20));
  drc_bufs26765 : INVD5BWP7T port map(I => n_1708, ZN => calc_buf_out(4));
  drc_bufs26771 : INVD5BWP7T port map(I => n_1714, ZN => calc_buf_out(19));
  drc_bufs26777 : INVD5BWP7T port map(I => n_1720, ZN => framebuffer_buf(15));
  drc_bufs26783 : INVD5BWP7T port map(I => n_1726, ZN => calc_buf_out(10));
  drc_bufs26789 : INVD5BWP7T port map(I => n_1732, ZN => calc_buf_out(5));
  drc_bufs26795 : INVD5BWP7T port map(I => n_1738, ZN => calc_buf_out(14));
  drc_bufs26801 : INVD5BWP7T port map(I => n_1744, ZN => calc_buf_out(13));
  drc_bufs26807 : INVD5BWP7T port map(I => n_1750, ZN => calc_buf_out(12));
  drc_bufs26813 : INVD5BWP7T port map(I => n_1756, ZN => calc_buf_out(11));
  drc_bufs26819 : INVD5BWP7T port map(I => n_1762, ZN => calc_buf_out(23));
  drc_bufs26825 : INVD5BWP7T port map(I => n_1768, ZN => calc_buf_out(6));
  drc_bufs26831 : INVD5BWP7T port map(I => n_1774, ZN => calc_buf_out(0));
  drc_bufs26837 : INVD5BWP7T port map(I => n_1780, ZN => calc_buf_out(16));
  drc_bufs26843 : INVD5BWP7T port map(I => n_1786, ZN => calc_buf_out(1));
  drc_bufs26849 : INVD5BWP7T port map(I => n_1792, ZN => framebuffer_buf(0));
  drc_bufs26855 : INVD5BWP7T port map(I => n_1798, ZN => calc_buf_out(8));
  drc_bufs26861 : INVD5BWP7T port map(I => n_1804, ZN => framebuffer_buf(1));
  drc_bufs26867 : INVD5BWP7T port map(I => n_1810, ZN => calc_buf_out(17));
  drc_bufs26873 : INVD5BWP7T port map(I => n_1816, ZN => calc_buf_out(9));
  state_reg_0 : DFKCND1BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_13, D => n_312, Q => state(0), QN => n_15);
  state_reg_2 : DFD1BWP7T port map(CP => CTS_14, D => n_251, Q => state(2), QN => n_89);
  counter_reg_4 : DFKCND1BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_14, D => new_counter(4), Q => counter(4), QN => n_70);
  counter_reg_0 : DFKCND1BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_14, D => new_counter(0), Q => counter(0), QN => n_252);
  counter_reg_3 : DFKCND1BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_14, D => new_counter(3), Q => counter(3), QN => n_327);
  counter_reg_5 : DFKCND1BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_14, D => new_counter(5), Q => counter(5), QN => n_242);
  state_reg_3 : DFD1BWP7T port map(CP => CTS_13, D => n_352, Q => state(3), QN => n_319);
  state_reg_1 : DFKCND1BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_13, D => n_287, Q => state(1), QN => n_143);
  counter_reg_7 : DFKCND1BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_14, D => new_counter(7), Q => counter(7), QN => n_504);
  counter_reg_2 : DFKCND1BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_14, D => new_counter(2), Q => counter(2), QN => n_355);
  counter_reg_1 : DFKCND1BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_14, D => new_counter(1), Q => counter(1), QN => n_246);
  counter_reg_6 : DFKCND1BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_14, D => new_counter(6), Q => counter(6), QN => n_393);
  calc_buf_out_reg_2 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_498, Q => calc_buf_out_2_2873, QN => n_742);
  framebuffer_buf_reg_157 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_585, Q => FE_PHN148_framebuffer_buf_157_3052, QN => n_748);
  framebuffer_buf_reg_156 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_583, Q => framebuffer_buf_156_3051, QN => n_754);
  framebuffer_buf_reg_155 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_13, D => n_539, Q => FE_PHN189_framebuffer_buf_155_3050, QN => n_760);
  framebuffer_buf_reg_154 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_13, D => n_514, Q => framebuffer_buf_154_3049, QN => n_766);
  framebuffer_buf_reg_153 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_608, Q => framebuffer_buf_153_3048, QN => n_772);
  framebuffer_buf_reg_152 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_614, Q => framebuffer_buf_152_3047, QN => n_778);
  framebuffer_buf_reg_151 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_623, Q => framebuffer_buf_151_3046, QN => n_784);
  framebuffer_buf_reg_150 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_580, Q => framebuffer_buf_150_3045, QN => n_790);
  framebuffer_buf_reg_149 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_584, Q => FE_PHN125_framebuffer_buf_149_3044, QN => n_796);
  framebuffer_buf_reg_148 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_586, Q => framebuffer_buf_148_3043, QN => n_802);
  framebuffer_buf_reg_147 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_537, Q => framebuffer_buf_147_3042, QN => n_808);
  framebuffer_buf_reg_146 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_538, Q => framebuffer_buf_146_3041, QN => n_814);
  framebuffer_buf_reg_145 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_523, Q => framebuffer_buf_145_3040, QN => n_820);
  framebuffer_buf_reg_144 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_524, Q => framebuffer_buf_144_3039, QN => n_826);
  framebuffer_buf_reg_143 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_525, Q => framebuffer_buf_143_3038, QN => n_832);
  framebuffer_buf_reg_142 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_526, Q => framebuffer_buf_142_3037, QN => n_838);
  framebuffer_buf_reg_141 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_510, Q => framebuffer_buf_141_3036, QN => n_844);
  framebuffer_buf_reg_140 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_511, Q => framebuffer_buf_140_3035, QN => n_850);
  framebuffer_buf_reg_139 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_657, Q => framebuffer_buf_139_3034, QN => n_856);
  framebuffer_buf_reg_138 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_660, Q => framebuffer_buf_138_3033, QN => n_862);
  calc_buf_out_reg_3 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_501, Q => calc_buf_out_3_2874, QN => n_868);
  framebuffer_buf_reg_136 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_640, Q => FE_PHN71_framebuffer_buf_136_3031, QN => n_874);
  framebuffer_buf_reg_135 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_579, Q => FE_PHN50_framebuffer_buf_135_3030, QN => n_880);
  framebuffer_buf_reg_134 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_662, Q => framebuffer_buf_134_3029, QN => n_886);
  framebuffer_buf_reg_133 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_588, Q => FE_PHN192_framebuffer_buf_133_3028, QN => n_892);
  framebuffer_buf_reg_132 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_591, Q => FE_PHN141_framebuffer_buf_132_3027, QN => n_898);
  framebuffer_buf_reg_131 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_593, Q => framebuffer_buf_131_3026, QN => n_904);
  framebuffer_buf_reg_130 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_598, Q => FE_PHN119_framebuffer_buf_130_3025, QN => n_910);
  calc_buf_out_reg_7 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_497, Q => calc_buf_out_7_2878, QN => n_916);
  framebuffer_buf_reg_128 : DFKCND0BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_13, D => n_639, Q => FE_PHN191_framebuffer_buf_128_3023, QN => n_922);
  framebuffer_buf_reg_127 : DFKCND0BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_13, D => n_620, Q => framebuffer_buf_127_3022, QN => n_928);
  framebuffer_buf_reg_126 : DFKCND0BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_13, D => n_621, Q => framebuffer_buf_126_3021, QN => n_934);
  framebuffer_buf_reg_125 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_622, Q => framebuffer_buf_125_3020, QN => n_940);
  framebuffer_buf_reg_124 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_14, D => n_629, Q => framebuffer_buf_124_3019, QN => n_946);
  framebuffer_buf_reg_123 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_550, Q => FE_PHN62_framebuffer_buf_123_3018, QN => n_952);
  framebuffer_buf_reg_122 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_551, Q => framebuffer_buf_122_3017, QN => n_958);
  calc_buf_out_reg_15 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_340, Q => calc_buf_out_15_2886, QN => n_964);
  framebuffer_buf_reg_120 : DFKCND0BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_13, D => n_545, Q => FE_PHN151_framebuffer_buf_120_3015, QN => n_970);
  framebuffer_buf_reg_119 : DFKCND0BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_13, D => n_546, Q => FE_PHN180_framebuffer_buf_119_3014, QN => n_976);
  framebuffer_buf_reg_118 : DFKCND0BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_13, D => n_547, Q => framebuffer_buf_118_3013, QN => n_982);
  framebuffer_buf_reg_115 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_515, Q => FE_PHN54_framebuffer_buf_115_3010, QN => n_988);
  framebuffer_buf_reg_114 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_516, Q => framebuffer_buf_114_3009, QN => n_994);
  framebuffer_buf_reg_113 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_512, Q => FE_PHN114_framebuffer_buf_113_3008, QN => n_1000);
  framebuffer_buf_reg_112 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_513, Q => framebuffer_buf_112_3007, QN => n_1006);
  framebuffer_buf_reg_7 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_385, Q => framebuffer_buf_7_2902, QN => n_1012);
  framebuffer_buf_reg_110 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_611, Q => framebuffer_buf_110_3005, QN => n_1018);
  framebuffer_buf_reg_109 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_568, Q => framebuffer_buf_109_3004, QN => n_1024);
  framebuffer_buf_reg_108 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_569, Q => framebuffer_buf_108_3003, QN => n_1030);
  framebuffer_buf_reg_107 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_13, D => n_570, Q => framebuffer_buf_107_3002, QN => n_1036);
  framebuffer_buf_reg_39 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_452, Q => framebuffer_buf_39_2934, QN => n_1042);
  framebuffer_buf_reg_103 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_506, Q => framebuffer_buf_103_2998, QN => n_1048);
  framebuffer_buf_reg_104 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_576, Q => framebuffer_buf_104_2999, QN => n_1054);
  framebuffer_buf_reg_40 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_451, Q => framebuffer_buf_40_2935, QN => n_1060);
  framebuffer_buf_reg_102 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_507, Q => framebuffer_buf_102_2997, QN => n_1066);
  framebuffer_buf_reg_101 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_646, Q => framebuffer_buf_101_2996, QN => n_1072);
  framebuffer_buf_reg_100 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_643, Q => framebuffer_buf_100_2995, QN => n_1078);
  framebuffer_buf_reg_99 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_647, Q => framebuffer_buf_99_2994, QN => n_1084);
  framebuffer_buf_reg_98 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_642, Q => framebuffer_buf_98_2993, QN => n_1090);
  framebuffer_buf_reg_97 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_565, Q => framebuffer_buf_97_2992, QN => n_1096);
  framebuffer_buf_reg_96 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_566, Q => framebuffer_buf_96_2991, QN => n_1102);
  framebuffer_buf_reg_95 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_552, Q => framebuffer_buf_95_2990, QN => n_1108);
  framebuffer_buf_reg_94 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_553, Q => framebuffer_buf_94_2989, QN => n_1114);
  framebuffer_buf_reg_93 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_555, Q => framebuffer_buf_93_2988, QN => n_1120);
  framebuffer_buf_reg_92 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_559, Q => framebuffer_buf_92_2987, QN => n_1126);
  framebuffer_buf_reg_91 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_607, Q => framebuffer_buf_91_2986, QN => n_1132);
  framebuffer_buf_reg_90 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_542, Q => framebuffer_buf_90_2985, QN => n_1138);
  framebuffer_buf_reg_89 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_527, Q => framebuffer_buf_89_2984, QN => n_1144);
  framebuffer_buf_reg_88 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_528, Q => framebuffer_buf_88_2983, QN => n_1150);
  framebuffer_buf_reg_87 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_529, Q => framebuffer_buf_87_2982, QN => n_1156);
  framebuffer_buf_reg_86 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_530, Q => framebuffer_buf_86_2981, QN => n_1162);
  framebuffer_buf_reg_85 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_554, Q => FE_PHN8_framebuffer_buf_85_2980, QN => n_1168);
  framebuffer_buf_reg_84 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_556, Q => framebuffer_buf_84_2979, QN => n_1174);
  framebuffer_buf_reg_83 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_557, Q => framebuffer_buf_83_2978, QN => n_1180);
  framebuffer_buf_reg_82 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_558, Q => framebuffer_buf_82_2977, QN => n_1186);
  framebuffer_buf_reg_81 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_562, Q => framebuffer_buf_81_2976, QN => n_1192);
  framebuffer_buf_reg_80 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_567, Q => framebuffer_buf_80_2975, QN => n_1198);
  framebuffer_buf_reg_105 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_575, Q => framebuffer_buf_105_3000, QN => n_1204);
  framebuffer_buf_reg_78 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_518, Q => framebuffer_buf_78_2973, QN => n_1210);
  framebuffer_buf_reg_77 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_604, Q => framebuffer_buf_77_2972, QN => n_1216);
  framebuffer_buf_reg_76 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_602, Q => framebuffer_buf_76_2971, QN => n_1222);
  framebuffer_buf_reg_106 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_13, D => n_571, Q => framebuffer_buf_106_3001, QN => n_1228);
  framebuffer_buf_reg_74 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_589, Q => framebuffer_buf_74_2969, QN => n_1234);
  framebuffer_buf_reg_73 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_533, Q => framebuffer_buf_73_2968, QN => n_1240);
  framebuffer_buf_reg_72 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_534, Q => framebuffer_buf_72_2967, QN => n_1246);
  framebuffer_buf_reg_8 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_423, Q => framebuffer_buf_8_2903, QN => n_1252);
  framebuffer_buf_reg_70 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_520, Q => framebuffer_buf_70_2965, QN => n_1258);
  framebuffer_buf_reg_69 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_521, Q => framebuffer_buf_69_2964, QN => n_1264);
  framebuffer_buf_reg_68 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_522, Q => framebuffer_buf_68_2963, QN => n_1270);
  framebuffer_buf_reg_67 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_508, Q => framebuffer_buf_67_2962, QN => n_1276);
  framebuffer_buf_reg_66 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_509, Q => framebuffer_buf_66_2961, QN => n_1282);
  framebuffer_buf_reg_65 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_649, Q => framebuffer_buf_65_2960, QN => n_1288);
  framebuffer_buf_reg_64 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_651, Q => framebuffer_buf_64_2959, QN => n_1294);
  framebuffer_buf_reg_63 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_655, Q => framebuffer_buf_63_2958, QN => n_1300);
  framebuffer_buf_reg_62 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_656, Q => framebuffer_buf_62_2957, QN => n_1306);
  framebuffer_buf_reg_61 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_628, Q => framebuffer_buf_61_2956, QN => n_1312);
  framebuffer_buf_reg_60 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_15, D => n_627, Q => framebuffer_buf_60_2955, QN => n_1318);
  framebuffer_buf_reg_59 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_599, Q => framebuffer_buf_59_2954, QN => n_1324);
  framebuffer_buf_reg_58 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_603, Q => FE_PHN87_framebuffer_buf_58_2953, QN => n_1330);
  framebuffer_buf_reg_57 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_605, Q => framebuffer_buf_57_2952, QN => n_1336);
  framebuffer_buf_reg_56 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_606, Q => framebuffer_buf_56_2951, QN => n_1342);
  framebuffer_buf_reg_137 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_661, Q => framebuffer_buf_137_3032, QN => n_1348);
  framebuffer_buf_reg_54 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_638, Q => framebuffer_buf_54_2949, QN => n_1354);
  framebuffer_buf_reg_53 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_615, Q => framebuffer_buf_53_2948, QN => n_1360);
  framebuffer_buf_reg_52 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_616, Q => framebuffer_buf_52_2947, QN => n_1366);
  framebuffer_buf_reg_129 : DFKCND0BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_13, D => n_636, Q => FE_PHN137_framebuffer_buf_129_3024, QN => n_1372);
  framebuffer_buf_reg_50 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_619, Q => framebuffer_buf_50_2945, QN => n_1378);
  framebuffer_buf_reg_49 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_474, Q => framebuffer_buf_49_2944, QN => n_1384);
  framebuffer_buf_reg_48 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_475, Q => framebuffer_buf_48_2943, QN => n_1390);
  framebuffer_buf_reg_121 : DFKCND0BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_13, D => n_544, Q => framebuffer_buf_121_3016, QN => n_1396);
  framebuffer_buf_reg_46 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_465, Q => framebuffer_buf_46_2941, QN => n_1402);
  framebuffer_buf_reg_45 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_466, Q => framebuffer_buf_45_2940, QN => n_1408);
  framebuffer_buf_reg_44 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_467, Q => framebuffer_buf_44_2939, QN => n_1414);
  framebuffer_buf_reg_41 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_478, Q => FE_PHN66_framebuffer_buf_41_2936, QN => n_1420);
  framebuffer_buf_reg_42 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_490, Q => framebuffer_buf_42_2937, QN => n_1426);
  framebuffer_buf_reg_9 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_438, Q => framebuffer_buf_9_2904, QN => n_1432);
  framebuffer_buf_reg_43 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_421, Q => framebuffer_buf_43_2938, QN => n_1438);
  framebuffer_buf_reg_111 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_617, Q => framebuffer_buf_111_3006, QN => n_1444);
  framebuffer_buf_reg_38 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_453, Q => framebuffer_buf_38_2933, QN => n_1450);
  framebuffer_buf_reg_37 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_424, Q => FE_PHN143_framebuffer_buf_37_2932, QN => n_1456);
  framebuffer_buf_reg_36 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_425, Q => framebuffer_buf_36_2931, QN => n_1462);
  framebuffer_buf_reg_35 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_426, Q => framebuffer_buf_35_2930, QN => n_1468);
  framebuffer_buf_reg_34 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_427, Q => framebuffer_buf_34_2929, QN => n_1474);
  framebuffer_buf_reg_33 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_430, Q => framebuffer_buf_33_2928, QN => n_1480);
  framebuffer_buf_reg_32 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_431, Q => framebuffer_buf_32_2927, QN => n_1486);
  framebuffer_buf_reg_31 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_445, Q => framebuffer_buf_31_2926, QN => n_1492);
  framebuffer_buf_reg_30 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_446, Q => framebuffer_buf_30_2925, QN => n_1498);
  framebuffer_buf_reg_29 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_439, Q => framebuffer_buf_29_2924, QN => n_1504);
  framebuffer_buf_reg_28 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_440, Q => FE_PHN69_framebuffer_buf_28_2923, QN => n_1510);
  framebuffer_buf_reg_79 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_517, Q => FE_PHN196_framebuffer_buf_79_2974, QN => n_1516);
  framebuffer_buf_reg_26 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_442, Q => framebuffer_buf_26_2921, QN => n_1522);
  framebuffer_buf_reg_75 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_594, Q => framebuffer_buf_75_2970, QN => n_1528);
  framebuffer_buf_reg_24 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_471, Q => framebuffer_buf_24_2919, QN => n_1534);
  framebuffer_buf_reg_71 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_519, Q => FE_PHN169_framebuffer_buf_71_2966, QN => n_1540);
  framebuffer_buf_reg_22 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_461, Q => framebuffer_buf_22_2917, QN => n_1546);
  framebuffer_buf_reg_21 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_462, Q => framebuffer_buf_21_2916, QN => n_1552);
  framebuffer_buf_reg_20 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_463, Q => framebuffer_buf_20_2915, QN => n_1558);
  framebuffer_buf_reg_19 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_456, Q => framebuffer_buf_19_2914, QN => n_1564);
  framebuffer_buf_reg_18 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_457, Q => framebuffer_buf_18_2913, QN => n_1570);
  framebuffer_buf_reg_17 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_447, Q => FE_PHN109_framebuffer_buf_17_2912, QN => n_1576);
  framebuffer_buf_reg_16 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_448, Q => framebuffer_buf_16_2911, QN => n_1582);
  framebuffer_buf_reg_55 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_633, Q => FE_PHN146_framebuffer_buf_55_2950, QN => n_1588);
  framebuffer_buf_reg_14 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_450, Q => framebuffer_buf_14_2909, QN => n_1594);
  framebuffer_buf_reg_51 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_618, Q => framebuffer_buf_51_2946, QN => n_1600);
  framebuffer_buf_reg_12 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_433, Q => framebuffer_buf_12_2907, QN => n_1606);
  framebuffer_buf_reg_10 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_437, Q => framebuffer_buf_10_2905, QN => n_1612);
  calc_buf_out_reg_18 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_354, Q => calc_buf_out_18_2889, QN => n_1618);
  framebuffer_buf_reg_11 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_434, Q => framebuffer_buf_11_2906, QN => n_1624);
  framebuffer_buf_reg_47 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_464, Q => framebuffer_buf_47_2942, QN => n_1630);
  framebuffer_buf_reg_13 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_432, Q => framebuffer_buf_13_2908, QN => n_1636);
  framebuffer_buf_reg_6 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_387, Q => framebuffer_buf_6_2901, QN => n_1642);
  framebuffer_buf_reg_5 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_392, Q => framebuffer_buf_5_2900, QN => n_1648);
  framebuffer_buf_reg_4 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_382, Q => framebuffer_buf_4_2899, QN => n_1654);
  framebuffer_buf_reg_3 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_383, Q => FE_PHN19_framebuffer_buf_3_2898, QN => n_1660);
  framebuffer_buf_reg_2 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_384, Q => framebuffer_buf_2_2897, QN => n_1666);
  framebuffer_buf_reg_27 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_441, Q => framebuffer_buf_27_2922, QN => n_1672);
  framebuffer_buf_reg_25 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_468, Q => framebuffer_buf_25_2920, QN => n_1678);
  framebuffer_buf_reg_23 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_14, D => n_479, Q => FE_PHN36_framebuffer_buf_23_2918, QN => n_1684);
  calc_buf_out_reg_22 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_339, Q => calc_buf_out_22_2893, QN => n_1690);
  calc_buf_out_reg_21 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_331, Q => calc_buf_out_21_2892, QN => n_1696);
  calc_buf_out_reg_20 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_332, Q => calc_buf_out_20_2891, QN => n_1702);
  calc_buf_out_reg_4 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_502, Q => calc_buf_out_4_2875, QN => n_1708);
  calc_buf_out_reg_19 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_330, Q => calc_buf_out_19_2890, QN => n_1714);
  framebuffer_buf_reg_15 : DFKCND0BWP7T port map(CN => FE_OFN3_n_0, CP => CTS_15, D => n_449, Q => framebuffer_buf_15_2910, QN => n_1720);
  calc_buf_out_reg_10 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_336, Q => FE_PHN68_calc_buf_out_10_2881, QN => n_1726);
  calc_buf_out_reg_5 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_492, Q => calc_buf_out_5_2876, QN => n_1732);
  calc_buf_out_reg_14 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_342, Q => calc_buf_out_14_2885, QN => n_1738);
  calc_buf_out_reg_13 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_351, Q => calc_buf_out_13_2884, QN => n_1744);
  calc_buf_out_reg_12 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_334, Q => calc_buf_out_12_2883, QN => n_1750);
  calc_buf_out_reg_11 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_335, Q => calc_buf_out_11_2882, QN => n_1756);
  calc_buf_out_reg_23 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_337, Q => calc_buf_out_23_2894, QN => n_1762);
  calc_buf_out_reg_6 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_496, Q => calc_buf_out_6_2877, QN => n_1768);
  calc_buf_out_reg_0 : DFKCND0BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_13, D => n_494, Q => calc_buf_out_0_2871, QN => n_1774);
  calc_buf_out_reg_16 : DFKCND0BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_13, D => n_344, Q => calc_buf_out_16_2887, QN => n_1780);
  calc_buf_out_reg_1 : DFKCND0BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_13, D => n_495, Q => calc_buf_out_1_2872, QN => n_1786);
  framebuffer_buf_reg_0 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_391, Q => framebuffer_buf_0_2895, QN => n_1792);
  calc_buf_out_reg_8 : DFKCND0BWP7T port map(CN => n_0, CP => CTS_13, D => n_348, Q => calc_buf_out_8_2879, QN => n_1798);
  framebuffer_buf_reg_1 : DFKCND0BWP7T port map(CN => FE_OFN1_n_0, CP => CTS_14, D => n_389, Q => framebuffer_buf_1_2896, QN => n_1804);
  calc_buf_out_reg_17 : DFKCND0BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_13, D => n_357, Q => calc_buf_out_17_2888, QN => n_1810);
  calc_buf_out_reg_9 : DFKCND0BWP7T port map(CN => FE_OFN2_n_0, CP => CTS_13, D => n_346, Q => FE_PHN16_calc_buf_out_9_2880, QN => n_1816);
  g27262 : INR2D1BWP7T port map(A1 => n_123, B1 => n_240, ZN => n_1820);
  g27263 : AO222D0BWP7T port map(A1 => n_379, A2 => counter(6), B1 => n_243, B2 => n_393, C1 => n_325, C2 => n_410, Z => n_1821);
  tie_0_cell : TIELBWP7T port map(ZN => FE_OFN4_framebuffer_buf_116);

end routed;
