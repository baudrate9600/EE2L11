library IEEE;
use IEEE.std_logic_1164.ALL;

entity mem_interface_tb is
end mem_interface_tb;

