configuration counter16_routed_cfg of counter16 is
   for routed
   end for;
end counter16_routed_cfg;
