
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture synthesised of memory is

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component LHQD1BWP7T
    port(E, D : in std_logic; Q : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCNQD1BWP7T
    port(CP, CN, D : in std_logic; Q : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component LNQD1BWP7T
    port(EN, D : in std_logic; Q : out std_logic);
  end component;

  component OAI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component CKND4BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component OAI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component LHD1BWP7T
    port(E, D : in std_logic; Q, QN : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component OAI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AOI211XD0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OAI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OA21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D4BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD4BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component DFD1BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CP, CN, D : in std_logic; Q, QN : out std_logic);
  end component;

  component DFKCND0BWP7T
    port(CP, CN, D : in std_logic; Q, QN : out std_logic);
  end component;

  signal new_row_buf : std_logic_vector(5 downto 0);
  signal new_counter : std_logic_vector(7 downto 0);
  signal counter : std_logic_vector(7 downto 0);
  signal row_buf : std_logic_vector(5 downto 0);
  signal state : std_logic_vector(3 downto 0);
  signal UNCONNECTED, UNCONNECTED0, UNCONNECTED1, UNCONNECTED2, UNCONNECTED3 : std_logic;
  signal UNCONNECTED4, UNCONNECTED5, UNCONNECTED6, calc_buf_out_0_2309, calc_buf_out_1_2310 : std_logic;
  signal calc_buf_out_2_2311, calc_buf_out_3_2312, calc_buf_out_4_2313, calc_buf_out_5_2314, calc_buf_out_6_2315 : std_logic;
  signal calc_buf_out_7_2316, calc_buf_out_8_2317, calc_buf_out_9_2318, calc_buf_out_10_2319, calc_buf_out_11_2320 : std_logic;
  signal calc_buf_out_12_2321, calc_buf_out_13_2322, calc_buf_out_14_2323, calc_buf_out_15_2324, calc_buf_out_16_2325 : std_logic;
  signal calc_buf_out_17_2326, calc_buf_out_18_2327, calc_buf_out_19_2328, calc_buf_out_20_2329, calc_buf_out_21_2330 : std_logic;
  signal calc_buf_out_22_2331, calc_buf_out_23_2332, framebuffer_buf_0_2333, framebuffer_buf_1_2334, framebuffer_buf_2_2335 : std_logic;
  signal framebuffer_buf_3_2336, framebuffer_buf_4_2337, framebuffer_buf_5_2338, framebuffer_buf_6_2339, framebuffer_buf_7_2340 : std_logic;
  signal framebuffer_buf_8_2341, framebuffer_buf_9_2342, framebuffer_buf_10_2343, framebuffer_buf_11_2344, framebuffer_buf_12_2345 : std_logic;
  signal framebuffer_buf_13_2346, framebuffer_buf_14_2347, framebuffer_buf_15_2348, framebuffer_buf_16_2349, framebuffer_buf_17_2350 : std_logic;
  signal framebuffer_buf_18_2351, framebuffer_buf_19_2352, framebuffer_buf_20_2353, framebuffer_buf_21_2354, framebuffer_buf_22_2355 : std_logic;
  signal framebuffer_buf_23_2356, framebuffer_buf_24_2357, framebuffer_buf_25_2358, framebuffer_buf_26_2359, framebuffer_buf_27_2360 : std_logic;
  signal framebuffer_buf_28_2361, framebuffer_buf_29_2362, framebuffer_buf_30_2363, framebuffer_buf_31_2364, framebuffer_buf_32_2365 : std_logic;
  signal framebuffer_buf_33_2366, framebuffer_buf_34_2367, framebuffer_buf_35_2368, framebuffer_buf_36_2369, framebuffer_buf_37_2370 : std_logic;
  signal framebuffer_buf_38_2371, framebuffer_buf_39_2372, framebuffer_buf_40_2373, framebuffer_buf_41_2374, framebuffer_buf_42_2375 : std_logic;
  signal framebuffer_buf_43_2376, framebuffer_buf_44_2377, framebuffer_buf_45_2378, framebuffer_buf_46_2379, framebuffer_buf_47_2380 : std_logic;
  signal framebuffer_buf_48_2381, framebuffer_buf_49_2382, framebuffer_buf_50_2383, framebuffer_buf_51_2384, framebuffer_buf_52_2385 : std_logic;
  signal framebuffer_buf_53_2386, framebuffer_buf_54_2387, framebuffer_buf_55_2388, framebuffer_buf_56_2389, framebuffer_buf_57_2390 : std_logic;
  signal framebuffer_buf_58_2391, framebuffer_buf_59_2392, framebuffer_buf_60_2393, framebuffer_buf_61_2394, framebuffer_buf_62_2395 : std_logic;
  signal framebuffer_buf_63_2396, framebuffer_buf_64_2397, framebuffer_buf_65_2398, framebuffer_buf_66_2399, framebuffer_buf_67_2400 : std_logic;
  signal framebuffer_buf_68_2401, framebuffer_buf_69_2402, framebuffer_buf_70_2403, framebuffer_buf_71_2404, framebuffer_buf_72_2405 : std_logic;
  signal framebuffer_buf_73_2406, framebuffer_buf_74_2407, framebuffer_buf_75_2408, framebuffer_buf_76_2409, framebuffer_buf_77_2410 : std_logic;
  signal framebuffer_buf_78_2411, framebuffer_buf_79_2412, framebuffer_buf_80_2413, framebuffer_buf_81_2414, framebuffer_buf_82_2415 : std_logic;
  signal framebuffer_buf_83_2416, framebuffer_buf_84_2417, framebuffer_buf_85_2418, framebuffer_buf_86_2419, framebuffer_buf_87_2420 : std_logic;
  signal framebuffer_buf_88_2421, framebuffer_buf_89_2422, framebuffer_buf_90_2423, framebuffer_buf_91_2424, framebuffer_buf_92_2425 : std_logic;
  signal framebuffer_buf_93_2426, framebuffer_buf_94_2427, framebuffer_buf_95_2428, framebuffer_buf_96_2429, framebuffer_buf_97_2430 : std_logic;
  signal framebuffer_buf_98_2431, framebuffer_buf_99_2432, framebuffer_buf_100_2433, framebuffer_buf_101_2434, framebuffer_buf_102_2435 : std_logic;
  signal framebuffer_buf_103_2436, framebuffer_buf_104_2437, framebuffer_buf_105_2438, framebuffer_buf_106_2439, framebuffer_buf_107_2440 : std_logic;
  signal framebuffer_buf_108_2441, framebuffer_buf_109_2442, framebuffer_buf_110_2443, framebuffer_buf_111_2444, framebuffer_buf_112_2445 : std_logic;
  signal framebuffer_buf_113_2446, framebuffer_buf_114_2447, framebuffer_buf_115_2448, framebuffer_buf_116_2449, framebuffer_buf_117_2450 : std_logic;
  signal framebuffer_buf_118_2451, framebuffer_buf_119_2452, framebuffer_buf_120_2453, framebuffer_buf_121_2454, framebuffer_buf_122_2455 : std_logic;
  signal framebuffer_buf_123_2456, framebuffer_buf_124_2457, framebuffer_buf_125_2458, framebuffer_buf_126_2459, framebuffer_buf_127_2460 : std_logic;
  signal framebuffer_buf_128_2461, framebuffer_buf_129_2462, framebuffer_buf_130_2463, framebuffer_buf_131_2464, framebuffer_buf_132_2465 : std_logic;
  signal framebuffer_buf_133_2466, framebuffer_buf_134_2467, framebuffer_buf_135_2468, framebuffer_buf_136_2469, framebuffer_buf_137_2470 : std_logic;
  signal framebuffer_buf_138_2471, framebuffer_buf_139_2472, framebuffer_buf_140_2473, framebuffer_buf_141_2474, framebuffer_buf_142_2475 : std_logic;
  signal framebuffer_buf_143_2476, framebuffer_buf_144_2477, framebuffer_buf_145_2478, framebuffer_buf_146_2479, framebuffer_buf_147_2480 : std_logic;
  signal framebuffer_buf_148_2481, framebuffer_buf_149_2482, framebuffer_buf_150_2483, framebuffer_buf_151_2484, framebuffer_buf_152_2485 : std_logic;
  signal framebuffer_buf_153_2486, framebuffer_buf_154_2487, framebuffer_buf_155_2488, framebuffer_buf_156_2489, framebuffer_buf_157_2490 : std_logic;
  signal n_0, n_1, n_2, n_4, n_5 : std_logic;
  signal n_6, n_7, n_8, n_9, n_12 : std_logic;
  signal n_13, n_14, n_15, n_16, n_17 : std_logic;
  signal n_18, n_21, n_22, n_23, n_25 : std_logic;
  signal n_26, n_27, n_29, n_30, n_31 : std_logic;
  signal n_32, n_33, n_34, n_35, n_36 : std_logic;
  signal n_44, n_45, n_46, n_49, n_52 : std_logic;
  signal n_53, n_54, n_55, n_56, n_58 : std_logic;
  signal n_59, n_60, n_61, n_62, n_63 : std_logic;
  signal n_65, n_67, n_68, n_69, n_70 : std_logic;
  signal n_71, n_72, n_74, n_75, n_76 : std_logic;
  signal n_77, n_78, n_79, n_80, n_81 : std_logic;
  signal n_82, n_83, n_84, n_85, n_86 : std_logic;
  signal n_88, n_90, n_91, n_92, n_93 : std_logic;
  signal n_94, n_95, n_96, n_97, n_98 : std_logic;
  signal n_99, n_100, n_101, n_102, n_103 : std_logic;
  signal n_104, n_105, n_106, n_107, n_109 : std_logic;
  signal n_110, n_111, n_112, n_113, n_114 : std_logic;
  signal n_115, n_116, n_117, n_118, n_119 : std_logic;
  signal n_120, n_121, n_122, n_123, n_124 : std_logic;
  signal n_125, n_126, n_127, n_128, n_129 : std_logic;
  signal n_130, n_131, n_132, n_133, n_134 : std_logic;
  signal n_135, n_136, n_137, n_138, n_139 : std_logic;
  signal n_140, n_141, n_142, n_143, n_144 : std_logic;
  signal n_145, n_146, n_147, n_148, n_149 : std_logic;
  signal n_150, n_151, n_152, n_153, n_154 : std_logic;
  signal n_155, n_156, n_157, n_158, n_159 : std_logic;
  signal n_160, n_161, n_162, n_170, n_173 : std_logic;
  signal n_174, n_175, n_176, n_177, n_178 : std_logic;
  signal n_179, n_180, n_181, n_182, n_183 : std_logic;
  signal n_184, n_186, n_187, n_188, n_189 : std_logic;
  signal n_190, n_191, n_192, n_193, n_194 : std_logic;
  signal n_195, n_196, n_197, n_198, n_199 : std_logic;
  signal n_200, n_201, n_202, n_203, n_204 : std_logic;
  signal n_205, n_206, n_207, n_208, n_209 : std_logic;
  signal n_210, n_211, n_212, n_213, n_214 : std_logic;
  signal n_215, n_216, n_217, n_218, n_219 : std_logic;
  signal n_220, n_221, n_222, n_223, n_224 : std_logic;
  signal n_225, n_226, n_227, n_228, n_229 : std_logic;
  signal n_230, n_231, n_232, n_233, n_234 : std_logic;
  signal n_235, n_236, n_237, n_238, n_239 : std_logic;
  signal n_240, n_241, n_242, n_243, n_244 : std_logic;
  signal n_245, n_246, n_247, n_248, n_249 : std_logic;
  signal n_250, n_251, n_252, n_253, n_254 : std_logic;
  signal n_255, n_256, n_257, n_258, n_259 : std_logic;
  signal n_260, n_261, n_262, n_263, n_264 : std_logic;
  signal n_265, n_266, n_267, n_268, n_269 : std_logic;
  signal n_270, n_271, n_272, n_273, n_274 : std_logic;
  signal n_275, n_276, n_277, n_278, n_279 : std_logic;
  signal n_280, n_281, n_282, n_283, n_284 : std_logic;
  signal n_285, n_286, n_287, n_288, n_289 : std_logic;
  signal n_290, n_291, n_292, n_293, n_294 : std_logic;
  signal n_295, n_296, n_297, n_298, n_299 : std_logic;
  signal n_300, n_301, n_302, n_303, n_304 : std_logic;
  signal n_305, n_306, n_307, n_308, n_309 : std_logic;
  signal n_310, n_311, n_312, n_313, n_314 : std_logic;
  signal n_315, n_316, n_317, n_318, n_319 : std_logic;
  signal n_320, n_321, n_322, n_323, n_324 : std_logic;
  signal n_325, n_326, n_327, n_328, n_329 : std_logic;
  signal n_330, n_331, n_332, n_333, n_334 : std_logic;
  signal n_335, n_336, n_337, n_338, n_339 : std_logic;
  signal n_340, n_341, n_342, n_343, n_344 : std_logic;
  signal n_345, n_346, n_347, n_348, n_349 : std_logic;
  signal n_350, n_351, n_352, n_353, n_354 : std_logic;
  signal n_355, n_356, n_357, n_358, n_359 : std_logic;
  signal n_360, n_361, n_362, n_363, n_364 : std_logic;
  signal n_365, n_366, n_367, n_368, n_369 : std_logic;
  signal n_370, n_371, n_372, n_373, n_374 : std_logic;
  signal n_375, n_376, n_377, n_378, n_379 : std_logic;
  signal n_380, n_381, n_382, n_383, n_384 : std_logic;
  signal n_385, n_386, n_387, n_388, n_389 : std_logic;
  signal n_390, n_391, n_392, n_393, n_394 : std_logic;
  signal n_395, n_396, n_397, n_398, n_399 : std_logic;
  signal n_400, n_401, n_402, n_403, n_404 : std_logic;
  signal n_405, n_406, n_407, n_408, n_409 : std_logic;
  signal n_410, n_411, n_412, n_413, n_414 : std_logic;
  signal n_415, n_416, n_417, n_418, n_419 : std_logic;
  signal n_420, n_421, n_422, n_423, n_424 : std_logic;
  signal n_425, n_426, n_427, n_428, n_429 : std_logic;
  signal n_430, n_431, n_432, n_433, n_434 : std_logic;
  signal n_435, n_436, n_437, n_438, n_439 : std_logic;
  signal n_443, n_444, n_445, n_446, n_459 : std_logic;
  signal n_460, n_461, n_462, n_463, n_465 : std_logic;
  signal n_466, n_467, n_468, n_469, n_470 : std_logic;
  signal n_471, n_472, n_493, n_496, n_502 : std_logic;
  signal n_508, n_514, n_520, n_526, n_532 : std_logic;
  signal n_538, n_544, n_550, n_556, n_562 : std_logic;
  signal n_568, n_574, n_580, n_586, n_592 : std_logic;
  signal n_598, n_604, n_610, n_616, n_622 : std_logic;
  signal n_628, n_634, n_640, n_646, n_652 : std_logic;
  signal n_658, n_664, n_670, n_676, n_682 : std_logic;
  signal n_688, n_694, n_700, n_706, n_712 : std_logic;
  signal n_718, n_724, n_730, n_736, n_742 : std_logic;
  signal n_748, n_754, n_760, n_766, n_772 : std_logic;
  signal n_778, n_784, n_790, n_796, n_802 : std_logic;
  signal n_808, n_814, n_820, n_826, n_832 : std_logic;
  signal n_838, n_844, n_850, n_856, n_862 : std_logic;
  signal n_868, n_874, n_880, n_886, n_892 : std_logic;
  signal n_898, n_904, n_910, n_916, n_922 : std_logic;
  signal n_928, n_934, n_940, n_946, n_952 : std_logic;
  signal n_958, n_964, n_970, n_976, n_982 : std_logic;
  signal n_988, n_994, n_1000, n_1006, n_1012 : std_logic;
  signal n_1018, n_1024, n_1030, n_1036, n_1042 : std_logic;
  signal n_1048, n_1054, n_1060, n_1066, n_1072 : std_logic;
  signal n_1078, n_1084, n_1090, n_1096, n_1102 : std_logic;
  signal n_1108, n_1114, n_1120, n_1126, n_1132 : std_logic;
  signal n_1138, n_1144, n_1150, n_1156, n_1162 : std_logic;
  signal n_1168, n_1174, n_1180, n_1186, n_1192 : std_logic;
  signal n_1198, n_1204, n_1210, n_1216, n_1222 : std_logic;
  signal n_1228, n_1234, n_1240, n_1246, n_1252 : std_logic;
  signal n_1258, n_1264, n_1270, n_1276, n_1282 : std_logic;
  signal n_1288, n_1294, n_1300, n_1306, n_1312 : std_logic;
  signal n_1318, n_1324, n_1330, n_1336, n_1342 : std_logic;
  signal n_1348, n_1354, n_1360, n_1366, n_1372 : std_logic;
  signal n_1378, n_1384, n_1390, n_1396, n_1402 : std_logic;
  signal n_1408, n_1414, n_1422, n_1428, n_1434 : std_logic;
  signal n_1440, n_1446, n_1452, n_1458, n_1464 : std_logic;
  signal n_1470, n_1476, n_1482, n_1488, n_1494 : std_logic;
  signal n_1500, n_1506, n_1512, n_1518, n_1524 : std_logic;
  signal n_1530, n_1536, n_1542, n_1548, n_1554 : std_logic;
  signal n_1560, n_1566, n_1572, n_1578, n_1584 : std_logic;
  signal n_1588, n_1589 : std_logic;

begin

  g23584 : AO22D0BWP7T port map(A1 => n_257, A2 => calc_buf_out_5_2314, B1 => sqi_data_in(5), B2 => n_461, Z => n_463);
  g23585 : AO22D0BWP7T port map(A1 => n_262, A2 => calc_buf_out_2_2311, B1 => sqi_data_in(2), B2 => n_461, Z => n_462);
  g23586 : AO22D0BWP7T port map(A1 => n_261, A2 => calc_buf_out_3_2312, B1 => sqi_data_in(3), B2 => n_461, Z => n_460);
  g23587 : AO22D0BWP7T port map(A1 => n_259, A2 => calc_buf_out_4_2313, B1 => sqi_data_in(4), B2 => n_461, Z => n_459);
  g23590 : AO22D0BWP7T port map(A1 => n_253, A2 => calc_buf_out_7_2316, B1 => sqi_data_in(7), B2 => n_461, Z => n_446);
  g23589 : AO22D0BWP7T port map(A1 => n_255, A2 => calc_buf_out_6_2315, B1 => sqi_data_in(6), B2 => n_461, Z => n_445);
  g23588 : AO22D0BWP7T port map(A1 => n_265, A2 => calc_buf_out_1_2310, B1 => sqi_data_in(1), B2 => n_461, Z => n_444);
  g23591 : AO22D0BWP7T port map(A1 => n_267, A2 => calc_buf_out_0_2309, B1 => sqi_data_in(0), B2 => n_461, Z => n_443);
  g23830 : MOAI22D0BWP7T port map(A1 => n_326, A2 => n_427, B1 => n_325, B2 => framebuffer_buf_84_2417, ZN => n_439);
  g23775 : MOAI22D0BWP7T port map(A1 => n_433, A2 => n_436, B1 => n_431, B2 => framebuffer_buf_117_2450, ZN => n_438);
  g23702 : MOAI22D0BWP7T port map(A1 => n_428, A2 => n_436, B1 => n_426, B2 => framebuffer_buf_133_2466, ZN => n_437);
  g23776 : MOAI22D0BWP7T port map(A1 => n_424, A2 => n_432, B1 => n_422, B2 => framebuffer_buf_14_2347, ZN => n_435);
  g23777 : MOAI22D0BWP7T port map(A1 => n_433, A2 => n_432, B1 => n_431, B2 => framebuffer_buf_118_2451, ZN => n_434);
  g23778 : MOAI22D0BWP7T port map(A1 => n_433, A2 => n_423, B1 => n_431, B2 => framebuffer_buf_119_2452, ZN => n_430);
  g23701 : MOAI22D0BWP7T port map(A1 => n_428, A2 => n_427, B1 => n_426, B2 => framebuffer_buf_132_2465, ZN => n_429);
  g23779 : MOAI22D0BWP7T port map(A1 => n_424, A2 => n_423, B1 => n_422, B2 => framebuffer_buf_15_2348, ZN => n_425);
  g23703 : MOAI22D0BWP7T port map(A1 => n_414, A2 => n_419, B1 => n_412, B2 => framebuffer_buf_136_2469, ZN => n_421);
  g23780 : MOAI22D0BWP7T port map(A1 => n_417, A2 => n_419, B1 => n_416, B2 => framebuffer_buf_120_2453, ZN => n_420);
  g23781 : MOAI22D0BWP7T port map(A1 => n_417, A2 => n_413, B1 => n_416, B2 => framebuffer_buf_121_2454, ZN => n_418);
  g23704 : MOAI22D0BWP7T port map(A1 => n_414, A2 => n_413, B1 => n_412, B2 => framebuffer_buf_137_2470, ZN => n_415);
  g23782 : MOAI22D0BWP7T port map(A1 => n_417, A2 => n_409, B1 => n_416, B2 => framebuffer_buf_122_2455, ZN => n_411);
  g23705 : MOAI22D0BWP7T port map(A1 => n_414, A2 => n_409, B1 => n_412, B2 => framebuffer_buf_138_2471, ZN => n_410);
  g23783 : MOAI22D0BWP7T port map(A1 => n_405, A2 => n_419, B1 => n_404, B2 => framebuffer_buf_16_2349, ZN => n_408);
  g23784 : MOAI22D0BWP7T port map(A1 => n_417, A2 => n_402, B1 => n_416, B2 => framebuffer_buf_123_2456, ZN => n_407);
  g23785 : MOAI22D0BWP7T port map(A1 => n_405, A2 => n_413, B1 => n_404, B2 => framebuffer_buf_17_2350, ZN => n_406);
  g23706 : MOAI22D0BWP7T port map(A1 => n_414, A2 => n_402, B1 => n_412, B2 => framebuffer_buf_139_2472, ZN => n_403);
  g23786 : MOAI22D0BWP7T port map(A1 => n_417, A2 => n_427, B1 => n_416, B2 => framebuffer_buf_124_2457, ZN => n_401);
  g23707 : MOAI22D0BWP7T port map(A1 => n_414, A2 => n_427, B1 => n_412, B2 => framebuffer_buf_140_2473, ZN => n_400);
  g23787 : MOAI22D0BWP7T port map(A1 => n_417, A2 => n_436, B1 => n_416, B2 => framebuffer_buf_125_2458, ZN => n_399);
  g23708 : MOAI22D0BWP7T port map(A1 => n_414, A2 => n_436, B1 => n_412, B2 => framebuffer_buf_141_2474, ZN => n_398);
  g23788 : MOAI22D0BWP7T port map(A1 => n_417, A2 => n_432, B1 => n_416, B2 => framebuffer_buf_126_2459, ZN => n_397);
  g23789 : MOAI22D0BWP7T port map(A1 => n_405, A2 => n_409, B1 => n_404, B2 => framebuffer_buf_18_2351, ZN => n_396);
  g23709 : MOAI22D0BWP7T port map(A1 => n_419, A2 => n_388, B1 => n_387, B2 => framebuffer_buf_56_2389, ZN => n_395);
  g23790 : MOAI22D0BWP7T port map(A1 => n_417, A2 => n_423, B1 => n_416, B2 => framebuffer_buf_127_2460, ZN => n_394);
  g23791 : MOAI22D0BWP7T port map(A1 => n_405, A2 => n_402, B1 => n_404, B2 => framebuffer_buf_19_2352, ZN => n_393);
  g23792 : MOAI22D0BWP7T port map(A1 => n_405, A2 => n_427, B1 => n_404, B2 => framebuffer_buf_20_2353, ZN => n_392);
  g23793 : MOAI22D0BWP7T port map(A1 => n_405, A2 => n_436, B1 => n_404, B2 => framebuffer_buf_21_2354, ZN => n_391);
  g23794 : MOAI22D0BWP7T port map(A1 => n_405, A2 => n_432, B1 => n_404, B2 => framebuffer_buf_22_2355, ZN => n_390);
  g23710 : MOAI22D0BWP7T port map(A1 => n_413, A2 => n_388, B1 => n_387, B2 => framebuffer_buf_57_2390, ZN => n_389);
  g23795 : MOAI22D0BWP7T port map(A1 => n_405, A2 => n_423, B1 => n_404, B2 => framebuffer_buf_23_2356, ZN => n_386);
  g23711 : MOAI22D0BWP7T port map(A1 => n_409, A2 => n_388, B1 => n_387, B2 => framebuffer_buf_58_2391, ZN => n_385);
  g23796 : MOAI22D0BWP7T port map(A1 => n_381, A2 => n_419, B1 => n_380, B2 => framebuffer_buf_144_2477, ZN => n_384);
  g23712 : MOAI22D0BWP7T port map(A1 => n_402, A2 => n_388, B1 => n_387, B2 => framebuffer_buf_59_2392, ZN => n_383);
  g23797 : MOAI22D0BWP7T port map(A1 => n_381, A2 => n_413, B1 => n_380, B2 => framebuffer_buf_145_2478, ZN => n_382);
  g23713 : MOAI22D0BWP7T port map(A1 => n_427, A2 => n_388, B1 => n_387, B2 => framebuffer_buf_60_2393, ZN => n_379);
  g23798 : MOAI22D0BWP7T port map(A1 => n_381, A2 => n_409, B1 => n_380, B2 => framebuffer_buf_146_2479, ZN => n_378);
  g23799 : MOAI22D0BWP7T port map(A1 => n_381, A2 => n_402, B1 => n_380, B2 => framebuffer_buf_147_2480, ZN => n_377);
  g23800 : MOAI22D0BWP7T port map(A1 => n_381, A2 => n_427, B1 => n_380, B2 => framebuffer_buf_148_2481, ZN => n_376);
  g23714 : MOAI22D0BWP7T port map(A1 => n_436, A2 => n_388, B1 => n_387, B2 => framebuffer_buf_61_2394, ZN => n_375);
  g23801 : MOAI22D0BWP7T port map(A1 => n_381, A2 => n_436, B1 => n_380, B2 => framebuffer_buf_149_2482, ZN => n_374);
  g23802 : MOAI22D0BWP7T port map(A1 => n_381, A2 => n_432, B1 => n_380, B2 => framebuffer_buf_150_2483, ZN => n_373);
  g23803 : MOAI22D0BWP7T port map(A1 => n_381, A2 => n_423, B1 => n_380, B2 => framebuffer_buf_151_2484, ZN => n_372);
  g23715 : MOAI22D0BWP7T port map(A1 => n_368, A2 => n_432, B1 => n_367, B2 => framebuffer_buf_110_2443, ZN => n_371);
  g23804 : MOAI22D0BWP7T port map(A1 => n_419, A2 => n_356, B1 => n_355, B2 => framebuffer_buf_32_2365, ZN => n_370);
  g23716 : MOAI22D0BWP7T port map(A1 => n_368, A2 => n_423, B1 => n_367, B2 => framebuffer_buf_111_2444, ZN => n_369);
  g23805 : MOAI22D0BWP7T port map(A1 => n_363, A2 => n_419, B1 => n_362, B2 => framebuffer_buf_152_2485, ZN => n_366);
  g23717 : MOAI22D0BWP7T port map(A1 => n_428, A2 => n_432, B1 => n_426, B2 => framebuffer_buf_134_2467, ZN => n_365);
  g23806 : MOAI22D0BWP7T port map(A1 => n_363, A2 => n_413, B1 => n_362, B2 => framebuffer_buf_153_2486, ZN => n_364);
  g23807 : MOAI22D0BWP7T port map(A1 => n_363, A2 => n_409, B1 => n_362, B2 => framebuffer_buf_154_2487, ZN => n_361);
  g23808 : MOAI22D0BWP7T port map(A1 => n_363, A2 => n_402, B1 => n_362, B2 => framebuffer_buf_155_2488, ZN => n_360);
  g23718 : MOAI22D0BWP7T port map(A1 => n_428, A2 => n_423, B1 => n_426, B2 => framebuffer_buf_135_2468, ZN => n_359);
  g23809 : MOAI22D0BWP7T port map(A1 => n_363, A2 => n_427, B1 => n_362, B2 => framebuffer_buf_156_2489, ZN => n_358);
  g23810 : MOAI22D0BWP7T port map(A1 => n_413, A2 => n_356, B1 => n_355, B2 => framebuffer_buf_33_2366, ZN => n_357);
  g23811 : MOAI22D0BWP7T port map(A1 => n_363, A2 => n_436, B1 => n_362, B2 => framebuffer_buf_157_2490, ZN => n_354);
  new_row_buf_reg_2 : LHQD1BWP7T port map(E => n_269, D => n_187, Q => new_row_buf(2));
  g23812 : MOAI22D0BWP7T port map(A1 => n_409, A2 => n_356, B1 => n_355, B2 => framebuffer_buf_34_2367, ZN => n_353);
  g23719 : MOAI22D0BWP7T port map(A1 => n_414, A2 => n_432, B1 => n_412, B2 => framebuffer_buf_142_2475, ZN => n_352);
  g23813 : MOAI22D0BWP7T port map(A1 => n_402, A2 => n_356, B1 => n_355, B2 => framebuffer_buf_35_2368, ZN => n_351);
  g23720 : MOAI22D0BWP7T port map(A1 => n_414, A2 => n_423, B1 => n_412, B2 => framebuffer_buf_143_2476, ZN => n_350);
  g23814 : MOAI22D0BWP7T port map(A1 => n_427, A2 => n_356, B1 => n_355, B2 => framebuffer_buf_36_2369, ZN => n_349);
  g23721 : MOAI22D0BWP7T port map(A1 => n_432, A2 => n_388, B1 => n_387, B2 => framebuffer_buf_62_2395, ZN => n_348);
  g23815 : MOAI22D0BWP7T port map(A1 => n_436, A2 => n_356, B1 => n_355, B2 => framebuffer_buf_37_2370, ZN => n_347);
  g23722 : MOAI22D0BWP7T port map(A1 => n_423, A2 => n_388, B1 => n_387, B2 => framebuffer_buf_63_2396, ZN => n_346);
  g23816 : MOAI22D0BWP7T port map(A1 => n_432, A2 => n_356, B1 => n_355, B2 => framebuffer_buf_38_2371, ZN => n_345);
  g23817 : MOAI22D0BWP7T port map(A1 => n_423, A2 => n_356, B1 => n_355, B2 => framebuffer_buf_39_2372, ZN => n_344);
  g23818 : MOAI22D0BWP7T port map(A1 => n_419, A2 => n_340, B1 => n_339, B2 => framebuffer_buf_48_2381, ZN => n_343);
  g23723 : MOAI22D0BWP7T port map(A1 => n_335, A2 => n_419, B1 => n_334, B2 => framebuffer_buf_72_2405, ZN => n_342);
  g23819 : MOAI22D0BWP7T port map(A1 => n_413, A2 => n_340, B1 => n_339, B2 => framebuffer_buf_49_2382, ZN => n_341);
  g23820 : MOAI22D0BWP7T port map(A1 => n_409, A2 => n_340, B1 => n_339, B2 => framebuffer_buf_50_2383, ZN => n_338);
  g23821 : MOAI22D0BWP7T port map(A1 => n_402, A2 => n_340, B1 => n_339, B2 => framebuffer_buf_51_2384, ZN => n_337);
  g23724 : MOAI22D0BWP7T port map(A1 => n_335, A2 => n_413, B1 => n_334, B2 => framebuffer_buf_73_2406, ZN => n_336);
  g23725 : MOAI22D0BWP7T port map(A1 => n_335, A2 => n_409, B1 => n_334, B2 => framebuffer_buf_74_2407, ZN => n_333);
  g23822 : MOAI22D0BWP7T port map(A1 => n_427, A2 => n_340, B1 => n_339, B2 => framebuffer_buf_52_2385, ZN => n_332);
  g23823 : MOAI22D0BWP7T port map(A1 => n_436, A2 => n_340, B1 => n_339, B2 => framebuffer_buf_53_2386, ZN => n_331);
  g23726 : MOAI22D0BWP7T port map(A1 => n_335, A2 => n_402, B1 => n_334, B2 => framebuffer_buf_75_2408, ZN => n_330);
  g23824 : MOAI22D0BWP7T port map(A1 => n_432, A2 => n_340, B1 => n_339, B2 => framebuffer_buf_54_2387, ZN => n_329);
  g23825 : MOAI22D0BWP7T port map(A1 => n_423, A2 => n_340, B1 => n_339, B2 => framebuffer_buf_55_2388, ZN => n_328);
  g23826 : MOAI22D0BWP7T port map(A1 => n_326, A2 => n_419, B1 => n_325, B2 => framebuffer_buf_80_2413, ZN => n_327);
  g23727 : MOAI22D0BWP7T port map(A1 => n_335, A2 => n_427, B1 => n_334, B2 => framebuffer_buf_76_2409, ZN => n_324);
  g23827 : MOAI22D0BWP7T port map(A1 => n_326, A2 => n_413, B1 => n_325, B2 => framebuffer_buf_81_2414, ZN => n_323);
  g23828 : MOAI22D0BWP7T port map(A1 => n_326, A2 => n_409, B1 => n_325, B2 => framebuffer_buf_82_2415, ZN => n_322);
  g23729 : MOAI22D0BWP7T port map(A1 => n_335, A2 => n_432, B1 => n_334, B2 => framebuffer_buf_78_2411, ZN => n_321);
  g23829 : MOAI22D0BWP7T port map(A1 => n_326, A2 => n_402, B1 => n_325, B2 => framebuffer_buf_83_2416, ZN => n_320);
  g23774 : MOAI22D0BWP7T port map(A1 => n_424, A2 => n_436, B1 => n_422, B2 => framebuffer_buf_13_2346, ZN => n_319);
  g23831 : MOAI22D0BWP7T port map(A1 => n_326, A2 => n_436, B1 => n_325, B2 => framebuffer_buf_85_2418, ZN => n_318);
  g23728 : MOAI22D0BWP7T port map(A1 => n_335, A2 => n_436, B1 => n_334, B2 => framebuffer_buf_77_2410, ZN => n_317);
  g23832 : MOAI22D0BWP7T port map(A1 => n_326, A2 => n_432, B1 => n_325, B2 => framebuffer_buf_86_2419, ZN => n_316);
  g23730 : MOAI22D0BWP7T port map(A1 => n_335, A2 => n_423, B1 => n_334, B2 => framebuffer_buf_79_2412, ZN => n_315);
  g23833 : MOAI22D0BWP7T port map(A1 => n_326, A2 => n_423, B1 => n_325, B2 => framebuffer_buf_87_2420, ZN => n_314);
  g23731 : MOAI22D0BWP7T port map(A1 => n_306, A2 => n_419, B1 => n_305, B2 => framebuffer_buf_64_2397, ZN => n_313);
  g23834 : MOAI22D0BWP7T port map(A1 => n_309, A2 => n_419, B1 => n_308, B2 => framebuffer_buf_88_2421, ZN => n_312);
  g23835 : MOAI22D0BWP7T port map(A1 => n_303, A2 => n_419, B1 => n_302, B2 => framebuffer_buf_0_2333, ZN => n_311);
  g23836 : MOAI22D0BWP7T port map(A1 => n_309, A2 => n_413, B1 => n_308, B2 => framebuffer_buf_89_2422, ZN => n_310);
  g23732 : MOAI22D0BWP7T port map(A1 => n_306, A2 => n_413, B1 => n_305, B2 => framebuffer_buf_65_2398, ZN => n_307);
  g23837 : MOAI22D0BWP7T port map(A1 => n_303, A2 => n_413, B1 => n_302, B2 => framebuffer_buf_1_2334, ZN => n_304);
  g23733 : MOAI22D0BWP7T port map(A1 => n_306, A2 => n_409, B1 => n_305, B2 => framebuffer_buf_66_2399, ZN => n_301);
  g23838 : MOAI22D0BWP7T port map(A1 => n_309, A2 => n_409, B1 => n_308, B2 => framebuffer_buf_90_2423, ZN => n_300);
  g23839 : MOAI22D0BWP7T port map(A1 => n_309, A2 => n_402, B1 => n_308, B2 => framebuffer_buf_91_2424, ZN => n_299);
  g23840 : MOAI22D0BWP7T port map(A1 => n_303, A2 => n_409, B1 => n_302, B2 => framebuffer_buf_2_2335, ZN => n_298);
  g23734 : MOAI22D0BWP7T port map(A1 => n_306, A2 => n_402, B1 => n_305, B2 => framebuffer_buf_67_2400, ZN => n_297);
  g23841 : MOAI22D0BWP7T port map(A1 => n_309, A2 => n_427, B1 => n_308, B2 => framebuffer_buf_92_2425, ZN => n_296);
  g23842 : MOAI22D0BWP7T port map(A1 => n_309, A2 => n_436, B1 => n_308, B2 => framebuffer_buf_93_2426, ZN => n_295);
  g23843 : MOAI22D0BWP7T port map(A1 => n_309, A2 => n_432, B1 => n_308, B2 => framebuffer_buf_94_2427, ZN => n_294);
  g23735 : MOAI22D0BWP7T port map(A1 => n_306, A2 => n_427, B1 => n_305, B2 => framebuffer_buf_68_2401, ZN => n_293);
  g23844 : MOAI22D0BWP7T port map(A1 => n_309, A2 => n_423, B1 => n_308, B2 => framebuffer_buf_95_2428, ZN => n_292);
  g23845 : MOAI22D0BWP7T port map(A1 => n_284, A2 => n_419, B1 => n_283, B2 => framebuffer_buf_96_2429, ZN => n_291);
  g23736 : MOAI22D0BWP7T port map(A1 => n_306, A2 => n_436, B1 => n_305, B2 => framebuffer_buf_69_2402, ZN => n_290);
  g23846 : MOAI22D0BWP7T port map(A1 => n_303, A2 => n_402, B1 => n_302, B2 => framebuffer_buf_3_2336, ZN => n_289);
  g23737 : MOAI22D0BWP7T port map(A1 => n_306, A2 => n_432, B1 => n_305, B2 => framebuffer_buf_70_2403, ZN => n_288);
  g23847 : MOAI22D0BWP7T port map(A1 => n_303, A2 => n_427, B1 => n_302, B2 => framebuffer_buf_4_2337, ZN => n_287);
  g23738 : MOAI22D0BWP7T port map(A1 => n_306, A2 => n_423, B1 => n_305, B2 => framebuffer_buf_71_2404, ZN => n_286);
  g23848 : MOAI22D0BWP7T port map(A1 => n_284, A2 => n_413, B1 => n_283, B2 => framebuffer_buf_97_2430, ZN => n_285);
  g23739 : MOAI22D0BWP7T port map(A1 => n_419, A2 => n_280, B1 => n_279, B2 => framebuffer_buf_24_2357, ZN => n_282);
  g23740 : MOAI22D0BWP7T port map(A1 => n_413, A2 => n_280, B1 => n_279, B2 => framebuffer_buf_25_2358, ZN => n_281);
  g23741 : MOAI22D0BWP7T port map(A1 => n_409, A2 => n_280, B1 => n_279, B2 => framebuffer_buf_26_2359, ZN => n_278);
  g23747 : MOAI22D0BWP7T port map(A1 => n_409, A2 => n_274, B1 => n_273, B2 => framebuffer_buf_42_2375, ZN => n_277);
  g23742 : MOAI22D0BWP7T port map(A1 => n_402, A2 => n_280, B1 => n_279, B2 => framebuffer_buf_27_2360, ZN => n_276);
  g23746 : MOAI22D0BWP7T port map(A1 => n_413, A2 => n_274, B1 => n_273, B2 => framebuffer_buf_41_2374, ZN => n_275);
  g23743 : MOAI22D0BWP7T port map(A1 => n_427, A2 => n_280, B1 => n_279, B2 => framebuffer_buf_28_2361, ZN => n_272);
  g23744 : MOAI22D0BWP7T port map(A1 => n_436, A2 => n_280, B1 => n_279, B2 => framebuffer_buf_29_2362, ZN => n_271);
  g23745 : MOAI22D0BWP7T port map(A1 => n_419, A2 => n_274, B1 => n_273, B2 => framebuffer_buf_40_2373, ZN => n_270);
  new_row_buf_reg_0 : LHQD1BWP7T port map(E => n_269, D => n_189, Q => new_row_buf(0));
  new_row_buf_reg_1 : LHQD1BWP7T port map(E => n_269, D => n_194, Q => new_row_buf(1));
  new_row_buf_reg_3 : LHQD1BWP7T port map(E => n_269, D => n_186, Q => new_row_buf(3));
  new_row_buf_reg_4 : LHQD1BWP7T port map(E => n_269, D => n_193, Q => new_row_buf(4));
  new_row_buf_reg_5 : LHQD1BWP7T port map(E => n_269, D => n_190, Q => new_row_buf(5));
  g23773 : MOAI22D0BWP7T port map(A1 => n_433, A2 => n_427, B1 => n_431, B2 => framebuffer_buf_116_2449, ZN => n_268);
  g23683 : ND2D0BWP7T port map(A1 => n_198, A2 => n_264, ZN => n_267);
  g23748 : MOAI22D0BWP7T port map(A1 => n_402, A2 => n_274, B1 => n_273, B2 => framebuffer_buf_43_2376, ZN => n_266);
  g23684 : ND2D0BWP7T port map(A1 => n_197, A2 => n_264, ZN => n_265);
  g23749 : MOAI22D0BWP7T port map(A1 => n_427, A2 => n_274, B1 => n_273, B2 => framebuffer_buf_44_2377, ZN => n_263);
  g23685 : ND2D0BWP7T port map(A1 => n_196, A2 => n_264, ZN => n_262);
  g23686 : ND2D0BWP7T port map(A1 => n_203, A2 => n_264, ZN => n_261);
  g23750 : MOAI22D0BWP7T port map(A1 => n_436, A2 => n_274, B1 => n_273, B2 => framebuffer_buf_45_2378, ZN => n_260);
  g23687 : ND2D0BWP7T port map(A1 => n_188, A2 => n_264, ZN => n_259);
  g23751 : MOAI22D0BWP7T port map(A1 => n_432, A2 => n_280, B1 => n_279, B2 => framebuffer_buf_30_2363, ZN => n_258);
  g23688 : ND2D0BWP7T port map(A1 => n_202, A2 => n_264, ZN => n_257);
  g23752 : MOAI22D0BWP7T port map(A1 => n_423, A2 => n_280, B1 => n_279, B2 => framebuffer_buf_31_2364, ZN => n_256);
  g23689 : ND2D0BWP7T port map(A1 => n_195, A2 => n_264, ZN => n_255);
  g23753 : MOAI22D0BWP7T port map(A1 => n_432, A2 => n_274, B1 => n_273, B2 => framebuffer_buf_46_2379, ZN => n_254);
  g23690 : ND2D0BWP7T port map(A1 => n_199, A2 => n_264, ZN => n_253);
  g23754 : MOAI22D0BWP7T port map(A1 => n_423, A2 => n_274, B1 => n_273, B2 => framebuffer_buf_47_2380, ZN => n_252);
  g23691 : MOAI22D0BWP7T port map(A1 => n_368, A2 => n_419, B1 => n_367, B2 => framebuffer_buf_104_2437, ZN => n_251);
  g23755 : MOAI22D0BWP7T port map(A1 => n_284, A2 => n_409, B1 => n_283, B2 => framebuffer_buf_98_2431, ZN => n_250);
  g23756 : MOAI22D0BWP7T port map(A1 => n_284, A2 => n_402, B1 => n_283, B2 => framebuffer_buf_99_2432, ZN => n_249);
  g23692 : MOAI22D0BWP7T port map(A1 => n_368, A2 => n_413, B1 => n_367, B2 => framebuffer_buf_105_2438, ZN => n_248);
  g23757 : MOAI22D0BWP7T port map(A1 => n_284, A2 => n_427, B1 => n_283, B2 => framebuffer_buf_100_2433, ZN => n_247);
  g23758 : MOAI22D0BWP7T port map(A1 => n_303, A2 => n_436, B1 => n_302, B2 => framebuffer_buf_5_2338, ZN => n_246);
  g23693 : MOAI22D0BWP7T port map(A1 => n_368, A2 => n_409, B1 => n_367, B2 => framebuffer_buf_106_2439, ZN => n_245);
  g23759 : MOAI22D0BWP7T port map(A1 => n_284, A2 => n_436, B1 => n_283, B2 => framebuffer_buf_101_2434, ZN => n_244);
  g23760 : MOAI22D0BWP7T port map(A1 => n_303, A2 => n_432, B1 => n_302, B2 => framebuffer_buf_6_2339, ZN => n_243);
  g23694 : MOAI22D0BWP7T port map(A1 => n_368, A2 => n_402, B1 => n_367, B2 => framebuffer_buf_107_2440, ZN => n_242);
  g23761 : MOAI22D0BWP7T port map(A1 => n_284, A2 => n_432, B1 => n_283, B2 => framebuffer_buf_102_2435, ZN => n_241);
  g23762 : MOAI22D0BWP7T port map(A1 => n_284, A2 => n_423, B1 => n_283, B2 => framebuffer_buf_103_2436, ZN => n_240);
  g23695 : MOAI22D0BWP7T port map(A1 => n_368, A2 => n_427, B1 => n_367, B2 => framebuffer_buf_108_2441, ZN => n_239);
  g23763 : MOAI22D0BWP7T port map(A1 => n_303, A2 => n_423, B1 => n_302, B2 => framebuffer_buf_7_2340, ZN => n_238);
  g23764 : MOAI22D0BWP7T port map(A1 => n_424, A2 => n_419, B1 => n_422, B2 => framebuffer_buf_8_2341, ZN => n_237);
  g23697 : MOAI22D0BWP7T port map(A1 => n_428, A2 => n_419, B1 => n_426, B2 => framebuffer_buf_128_2461, ZN => n_236);
  g23765 : MOAI22D0BWP7T port map(A1 => n_424, A2 => n_413, B1 => n_422, B2 => framebuffer_buf_9_2342, ZN => n_235);
  g23766 : MOAI22D0BWP7T port map(A1 => n_424, A2 => n_409, B1 => n_422, B2 => framebuffer_buf_10_2343, ZN => n_234);
  g23767 : MOAI22D0BWP7T port map(A1 => n_433, A2 => n_419, B1 => n_431, B2 => framebuffer_buf_112_2445, ZN => n_233);
  g23696 : MOAI22D0BWP7T port map(A1 => n_368, A2 => n_436, B1 => n_367, B2 => framebuffer_buf_109_2442, ZN => n_232);
  g23768 : MOAI22D0BWP7T port map(A1 => n_424, A2 => n_402, B1 => n_422, B2 => framebuffer_buf_11_2344, ZN => n_231);
  g23698 : MOAI22D0BWP7T port map(A1 => n_428, A2 => n_413, B1 => n_426, B2 => framebuffer_buf_129_2462, ZN => n_230);
  g23769 : MOAI22D0BWP7T port map(A1 => n_433, A2 => n_413, B1 => n_431, B2 => framebuffer_buf_113_2446, ZN => n_229);
  g23699 : MOAI22D0BWP7T port map(A1 => n_428, A2 => n_409, B1 => n_426, B2 => framebuffer_buf_130_2463, ZN => n_228);
  g23770 : MOAI22D0BWP7T port map(A1 => n_433, A2 => n_409, B1 => n_431, B2 => framebuffer_buf_114_2447, ZN => n_227);
  g23771 : MOAI22D0BWP7T port map(A1 => n_424, A2 => n_427, B1 => n_422, B2 => framebuffer_buf_12_2345, ZN => n_226);
  g23772 : MOAI22D0BWP7T port map(A1 => n_433, A2 => n_402, B1 => n_431, B2 => framebuffer_buf_115_2448, ZN => n_225);
  g23700 : MOAI22D0BWP7T port map(A1 => n_428, A2 => n_402, B1 => n_426, B2 => framebuffer_buf_131_2464, ZN => n_224);
  counter_reg_7 : DFKCNQD1BWP7T port map(CP => clk, CN => n_2, D => new_counter(7), Q => counter(7));
  g23865 : AO22D0BWP7T port map(A1 => n_221, A2 => calc_buf_out_9_2318, B1 => sqi_data_in(1), B2 => n_220, Z => n_223);
  g23869 : AO22D0BWP7T port map(A1 => n_221, A2 => calc_buf_out_13_2322, B1 => sqi_data_in(5), B2 => n_220, Z => n_222);
  g23867 : AO22D0BWP7T port map(A1 => n_221, A2 => calc_buf_out_11_2320, B1 => sqi_data_in(3), B2 => n_220, Z => n_219);
  g23864 : AO22D0BWP7T port map(A1 => n_212, A2 => calc_buf_out_23_2332, B1 => sqi_data_in(7), B2 => n_211, Z => n_218);
  g23871 : AO22D0BWP7T port map(A1 => n_221, A2 => calc_buf_out_14_2323, B1 => sqi_data_in(6), B2 => n_220, Z => n_217);
  g23866 : AO22D0BWP7T port map(A1 => n_221, A2 => calc_buf_out_10_2319, B1 => sqi_data_in(2), B2 => n_220, Z => n_216);
  g23868 : AO22D0BWP7T port map(A1 => n_221, A2 => calc_buf_out_12_2321, B1 => sqi_data_in(4), B2 => n_220, Z => n_215);
  g23870 : AO22D0BWP7T port map(A1 => n_221, A2 => calc_buf_out_15_2324, B1 => sqi_data_in(7), B2 => n_220, Z => n_214);
  g23876 : AO22D0BWP7T port map(A1 => n_212, A2 => calc_buf_out_20_2329, B1 => sqi_data_in(4), B2 => n_211, Z => n_213);
  g23873 : AO22D0BWP7T port map(A1 => n_212, A2 => calc_buf_out_17_2326, B1 => sqi_data_in(1), B2 => n_211, Z => n_210);
  g23874 : AO22D0BWP7T port map(A1 => n_212, A2 => calc_buf_out_18_2327, B1 => sqi_data_in(2), B2 => n_211, Z => n_209);
  g23875 : AO22D0BWP7T port map(A1 => n_212, A2 => calc_buf_out_19_2328, B1 => sqi_data_in(3), B2 => n_211, Z => n_208);
  g23872 : AO22D0BWP7T port map(A1 => n_212, A2 => calc_buf_out_16_2325, B1 => sqi_data_in(0), B2 => n_211, Z => n_207);
  g23877 : AO22D0BWP7T port map(A1 => n_212, A2 => calc_buf_out_21_2330, B1 => sqi_data_in(5), B2 => n_211, Z => n_206);
  g23878 : AO22D0BWP7T port map(A1 => n_212, A2 => calc_buf_out_22_2331, B1 => sqi_data_in(6), B2 => n_211, Z => n_205);
  g23879 : AO22D0BWP7T port map(A1 => n_221, A2 => calc_buf_out_8_2317, B1 => sqi_data_in(0), B2 => n_220, Z => n_204);
  g23861 : OAI31D0BWP7T port map(A1 => sqi_data_in(3), A2 => n_303, A3 => n_201, B => n_200, ZN => n_203);
  g23856 : OAI31D0BWP7T port map(A1 => sqi_data_in(5), A2 => n_303, A3 => n_201, B => n_200, ZN => n_202);
  g23857 : OAI31D0BWP7T port map(A1 => sqi_data_in(7), A2 => n_303, A3 => n_201, B => n_200, ZN => n_199);
  g23858 : OAI31D0BWP7T port map(A1 => sqi_data_in(0), A2 => n_303, A3 => n_201, B => n_200, ZN => n_198);
  g23859 : OAI31D0BWP7T port map(A1 => sqi_data_in(1), A2 => n_303, A3 => n_201, B => n_200, ZN => n_197);
  g23860 : OAI31D0BWP7T port map(A1 => sqi_data_in(2), A2 => n_303, A3 => n_201, B => n_200, ZN => n_196);
  g23849 : OAI31D0BWP7T port map(A1 => sqi_data_in(6), A2 => n_303, A3 => n_201, B => n_200, ZN => n_195);
  g23899 : AO22D0BWP7T port map(A1 => n_192, A2 => row_buf(1), B1 => sqi_data_in(1), B2 => n_191, Z => n_194);
  g23902 : AO22D0BWP7T port map(A1 => n_192, A2 => row_buf(4), B1 => sqi_data_in(4), B2 => n_191, Z => n_193);
  g23897 : AO22D0BWP7T port map(A1 => n_192, A2 => row_buf(5), B1 => sqi_data_in(5), B2 => n_191, Z => n_190);
  g23898 : AO22D0BWP7T port map(A1 => n_192, A2 => row_buf(0), B1 => sqi_data_in(0), B2 => n_191, Z => n_189);
  g23862 : OAI31D0BWP7T port map(A1 => sqi_data_in(4), A2 => n_303, A3 => n_201, B => n_200, ZN => n_188);
  g23900 : AO22D0BWP7T port map(A1 => n_192, A2 => row_buf(2), B1 => sqi_data_in(2), B2 => n_191, Z => n_187);
  g23901 : AO22D0BWP7T port map(A1 => n_192, A2 => row_buf(3), B1 => sqi_data_in(3), B2 => n_191, Z => n_186);
  g23892 : OAI21D0BWP7T port map(A1 => n_84, A2 => n_184, B => n_183, ZN => n_305);
  g23886 : OAI21D0BWP7T port map(A1 => n_75, A2 => n_184, B => n_183, ZN => n_279);
  g23887 : OAI21D0BWP7T port map(A1 => n_82, A2 => n_184, B => n_183, ZN => n_367);
  g23888 : OAI21D0BWP7T port map(A1 => n_111, A2 => n_184, B => n_183, ZN => n_426);
  g23889 : OAI21D0BWP7T port map(A1 => n_91, A2 => n_184, B => n_183, ZN => n_412);
  g23890 : OAI21D0BWP7T port map(A1 => n_77, A2 => n_184, B => n_183, ZN => n_387);
  g23891 : OAI21D0BWP7T port map(A1 => n_60, A2 => n_184, B => n_183, ZN => n_334);
  state_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => n_2, D => n_173, Q => state(0));
  new_counter_reg_7 : LNQD1BWP7T port map(EN => n_176, D => n_177, Q => new_counter(7));
  g23903 : OAI21D0BWP7T port map(A1 => n_95, A2 => n_184, B => n_183, ZN => n_362);
  state_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => n_2, D => n_174, Q => state(1));
  g23904 : OAI21D0BWP7T port map(A1 => n_112, A2 => n_184, B => n_183, ZN => n_380);
  g23905 : OAI21D0BWP7T port map(A1 => n_76, A2 => n_184, B => n_183, ZN => n_339);
  g23906 : OAI21D0BWP7T port map(A1 => n_182, A2 => n_184, B => n_183, ZN => n_404);
  g23907 : OAI21D0BWP7T port map(A1 => n_79, A2 => n_184, B => n_183, ZN => n_325);
  g23893 : OAI21D0BWP7T port map(A1 => n_83, A2 => n_184, B => n_183, ZN => n_273);
  g23909 : OAI21D0BWP7T port map(A1 => n_86, A2 => n_184, B => n_183, ZN => n_431);
  g23910 : OAI21D0BWP7T port map(A1 => n_92, A2 => n_184, B => n_183, ZN => n_416);
  g23911 : OAI21D0BWP7T port map(A1 => n_81, A2 => n_184, B => n_183, ZN => n_355);
  g23912 : OAI21D0BWP7T port map(A1 => n_68, A2 => n_184, B => n_183, ZN => n_283);
  g23913 : OAI21D0BWP7T port map(A1 => n_180, A2 => n_184, B => n_183, ZN => n_422);
  g23914 : OAI21D0BWP7T port map(A1 => n_80, A2 => n_184, B => n_183, ZN => n_302);
  g23908 : OAI21D0BWP7T port map(A1 => n_85, A2 => n_184, B => n_183, ZN => n_308);
  g23918 : OAI211D1BWP7T port map(A1 => n_181, A2 => n_182, B => n_179, C => n_178, ZN => n_212);
  g23919 : OAI211D1BWP7T port map(A1 => n_181, A2 => n_180, B => n_179, C => n_178, ZN => n_221);
  g23952 : AO21D0BWP7T port map(A1 => n_154, A2 => counter(7), B => n_139, Z => n_177);
  g23917 : ND2D1BWP7T port map(A1 => n_179, A2 => n_181, ZN => n_200);
  new_counter_reg_6 : LNQD1BWP7T port map(EN => n_176, D => n_170, Q => new_counter(6));
  g23933 : OR2D0BWP7T port map(A1 => n_175, A2 => n_155, Z => n_192);
  g23920 : NR3D0BWP7T port map(A1 => n_175, A2 => n_65, A3 => n_191, ZN => n_183);
  new_counter_reg_3 : LNQD1BWP7T port map(EN => n_176, D => n_162, Q => new_counter(3));
  g23915 : ND4D0BWP7T port map(A1 => n_143, A2 => n_146, A3 => n_148, A4 => n_61, ZN => n_174);
  new_counter_reg_0 : LNQD1BWP7T port map(EN => n_176, D => n_145, Q => new_counter(0));
  new_counter_reg_1 : LNQD1BWP7T port map(EN => n_176, D => n_160, Q => new_counter(1));
  new_counter_reg_5 : LNQD1BWP7T port map(EN => n_176, D => n_156, Q => new_counter(5));
  g23931 : IND4D0BWP7T port map(A1 => n_147, B1 => n_93, B2 => n_150, B3 => n_151, ZN => n_173);
  new_counter_reg_2 : LNQD1BWP7T port map(EN => n_176, D => n_159, Q => new_counter(2));
  new_counter_reg_4 : LNQD1BWP7T port map(EN => n_176, D => n_157, Q => new_counter(4));
  g23927 : INVD1BWP7T port map(I => n_179, ZN => n_201);
  g23951 : CKND4BWP7T port map(I => n_465, ZN => sqi_data_out(7));
  g23949 : CKND4BWP7T port map(I => n_466, ZN => sqi_data_out(0));
  g23962 : OAI32D0BWP7T port map(A1 => counter(6), A2 => n_161, A3 => n_138, B1 => n_137, B2 => n_153, ZN => n_170);
  g23953 : IND2D1BWP7T port map(A1 => n_1588, B1 => n_178, ZN => n_175);
  g23934 : NR3D0BWP7T port map(A1 => n_1588, A2 => n_31, A3 => n_191, ZN => n_179);
  g23936 : CKND4BWP7T port map(I => n_472, ZN => sqi_data_out(2));
  g23938 : CKND4BWP7T port map(I => n_471, ZN => sqi_data_out(3));
  g23940 : CKND4BWP7T port map(I => n_470, ZN => sqi_data_out(4));
  g23942 : CKND4BWP7T port map(I => n_469, ZN => sqi_data_out(1));
  g23944 : CKND4BWP7T port map(I => n_468, ZN => sqi_data_out(5));
  g23946 : CKND4BWP7T port map(I => n_467, ZN => sqi_data_out(6));
  g23961 : OAI32D0BWP7T port map(A1 => counter(3), A2 => n_114, A3 => n_161, B1 => n_32, B2 => n_115, ZN => n_162);
  sqi_data_out_reg_7 : LHD1BWP7T port map(E => n_158, D => n_90, Q => UNCONNECTED, QN => n_465);
  g23965 : OAI32D0BWP7T port map(A1 => counter(1), A2 => n_144, A3 => n_161, B1 => n_96, B2 => n_116, ZN => n_160);
  g23958 : OAI32D0BWP7T port map(A1 => counter(2), A2 => n_122, A3 => n_161, B1 => n_16, B2 => n_123, ZN => n_159);
  sqi_data_out_reg_0 : LHD1BWP7T port map(E => n_158, D => n_113, Q => UNCONNECTED0, QN => n_466);
  g23963 : OAI32D0BWP7T port map(A1 => counter(4), A2 => n_119, A3 => n_161, B1 => n_15, B2 => n_120, ZN => n_157);
  g23964 : OAI32D0BWP7T port map(A1 => counter(5), A2 => n_117, A3 => n_161, B1 => n_22, B2 => n_118, ZN => n_156);
  g23955 : NR2D0BWP7T port map(A1 => n_142, A2 => n_155, ZN => n_176);
  sqi_data_out_reg_6 : LHD1BWP7T port map(E => n_158, D => n_128, Q => UNCONNECTED1, QN => n_467);
  g23969 : OAI21D0BWP7T port map(A1 => n_94, A2 => counter(6), B => n_153, ZN => n_154);
  g23932 : ND4D0BWP7T port map(A1 => n_125, A2 => n_151, A3 => n_141, A4 => n_2, ZN => n_152);
  sqi_data_out_reg_2 : LHD1BWP7T port map(E => n_158, D => n_140, Q => UNCONNECTED2, QN => n_472);
  sqi_data_out_reg_3 : LHD1BWP7T port map(E => n_158, D => n_131, Q => UNCONNECTED3, QN => n_471);
  sqi_data_out_reg_4 : LHD1BWP7T port map(E => n_158, D => n_129, Q => UNCONNECTED4, QN => n_470);
  sqi_data_out_reg_1 : LHD1BWP7T port map(E => n_158, D => n_136, Q => UNCONNECTED5, QN => n_469);
  sqi_data_out_reg_5 : LHD1BWP7T port map(E => n_158, D => n_130, Q => UNCONNECTED6, QN => n_468);
  state_reg_2 : DFQD1BWP7T port map(CP => clk, D => n_127, Q => state(2));
  g23954 : ND4D0BWP7T port map(A1 => n_133, A2 => n_149, A3 => n_148, A4 => n_55, ZN => n_269);
  g23966 : OAI211D0BWP7T port map(A1 => sqi_finished, A2 => n_184, B => n_106, C => n_132, ZN => n_147);
  g23970 : AOI211XD0BWP7T port map(A1 => n_104, A2 => n_99, B => n_109, C => n_56, ZN => n_146);
  g23971 : OAI222D0BWP7T port map(A1 => n_110, A2 => n_178, B1 => n_144, B2 => n_107, C1 => counter(0), C2 => n_161, ZN => n_145);
  g23956 : AOI22D0BWP7T port map(A1 => n_124, A2 => n_46, B1 => n_105, B2 => n_45, ZN => n_143);
  g23957 : OAI211D0BWP7T port map(A1 => n_178, A2 => n_70, B => n_126, C => n_141, ZN => n_142);
  g23973 : AO22D0BWP7T port map(A1 => n_135, A2 => calc_buf_in(1), B1 => row_buf(2), B2 => n_134, Z => n_140);
  g23968 : NR4D0BWP7T port map(A1 => n_138, A2 => n_161, A3 => n_137, A4 => counter(7), ZN => n_139);
  g23972 : AO22D0BWP7T port map(A1 => n_135, A2 => calc_buf_in(0), B1 => row_buf(1), B2 => n_134, Z => n_136);
  g23960 : ND3D0BWP7T port map(A1 => n_133, A2 => n_149, A3 => n_132, ZN => n_158);
  g23974 : AO22D0BWP7T port map(A1 => n_135, A2 => calc_buf_in(2), B1 => row_buf(3), B2 => n_134, Z => n_131);
  g23975 : AO22D0BWP7T port map(A1 => n_135, A2 => calc_buf_in(4), B1 => row_buf(5), B2 => n_134, Z => n_130);
  g23976 : AO22D0BWP7T port map(A1 => n_135, A2 => calc_buf_in(3), B1 => row_buf(4), B2 => n_134, Z => n_129);
  g23977 : AO22D0BWP7T port map(A1 => n_135, A2 => calc_buf_in(5), B1 => calc_buf_in(0), B2 => n_134, Z => n_128);
  g23947 : ND4D0BWP7T port map(A1 => n_126, A2 => n_493, A3 => n_184, A4 => n_2, ZN => n_127);
  g23986 : AOI21D0BWP7T port map(A1 => n_138, A2 => n_155, B => n_121, ZN => n_153);
  g23967 : NR2D0BWP7T port map(A1 => n_124, A2 => n_103, ZN => n_125);
  g23978 : AOI21D0BWP7T port map(A1 => n_155, A2 => n_122, B => n_121, ZN => n_123);
  g23979 : AOI21D0BWP7T port map(A1 => n_155, A2 => n_119, B => n_121, ZN => n_120);
  g23984 : AOI21D0BWP7T port map(A1 => n_117, A2 => n_155, B => n_121, ZN => n_118);
  g23983 : AOI21D0BWP7T port map(A1 => n_155, A2 => n_144, B => n_121, ZN => n_116);
  g23982 : AOI21D0BWP7T port map(A1 => n_155, A2 => n_114, B => n_121, ZN => n_115);
  g24012 : INR2D0BWP7T port map(A1 => row_buf(0), B1 => n_149, ZN => n_113);
  g23980 : NR2D0BWP7T port map(A1 => n_88, A2 => n_155, ZN => n_133);
  g23989 : INVD1BWP7T port map(I => n_112, ZN => n_381);
  g23990 : INVD1BWP7T port map(I => n_111, ZN => n_428);
  g23992 : ND2D1BWP7T port map(A1 => n_110, A2 => n_69, ZN => n_264);
  g23999 : AOI22D0BWP7T port map(A1 => n_151, A2 => n_101, B1 => n_178, B2 => n_100, ZN => n_109);
  g23996 : INVD0BWP7T port map(I => n_121, ZN => n_107);
  g24001 : AOI22D0BWP7T port map(A1 => n_105, A2 => n_44, B1 => n_54, B2 => n_104, ZN => n_106);
  g24028 : NR2XD0BWP7T port map(A1 => n_405, A2 => n_181, ZN => n_211);
  g23998 : OAI222D0BWP7T port map(A1 => ce, A2 => n_102, B1 => n_101, B2 => n_100, C1 => n_99, C2 => n_35, ZN => n_103);
  g23985 : AOI22D0BWP7T port map(A1 => n_98, A2 => n_30, B1 => n_62, B2 => ce, ZN => n_126);
  g23981 : OAI21D0BWP7T port map(A1 => n_98, A2 => n_150, B => n_21, ZN => n_124);
  g23995 : NR2XD0BWP7T port map(A1 => n_97, A2 => counter(1), ZN => n_111);
  g23994 : NR2XD0BWP7T port map(A1 => n_97, A2 => n_96, ZN => n_112);
  g23987 : INVD1BWP7T port map(I => n_95, ZN => n_363);
  g24002 : OAI211D0BWP7T port map(A1 => sqi_finished, A2 => n_94, B => n_150, C => n_178, ZN => n_121);
  g24003 : ND3D0BWP7T port map(A1 => n_148, A2 => n_101, A3 => n_93, ZN => n_135);
  g24005 : INVD1BWP7T port map(I => n_92, ZN => n_417);
  g23988 : INVD1BWP7T port map(I => n_91, ZN => n_414);
  g24010 : INR2D0BWP7T port map(A1 => calc_buf_in(1), B1 => n_149, ZN => n_90);
  row_buf_reg_4 : DFKCNQD1BWP7T port map(CP => clk, CN => n_2, D => new_row_buf(4), Q => row_buf(4));
  g24024 : OA21D0BWP7T port map(A1 => n_101, A2 => n_36, B => n_148, Z => n_132);
  row_buf_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => n_2, D => new_row_buf(1), Q => row_buf(1));
  row_buf_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => n_2, D => new_row_buf(3), Q => row_buf(3));
  row_buf_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => n_2, D => new_row_buf(0), Q => row_buf(0));
  row_buf_reg_5 : DFKCNQD1BWP7T port map(CP => clk, CN => n_2, D => new_row_buf(5), Q => row_buf(5));
  row_buf_reg_2 : DFKCNQD1BWP7T port map(CP => clk, CN => n_2, D => new_row_buf(2), Q => row_buf(2));
  g24013 : IND2D0BWP7T port map(A1 => n_117, B1 => counter(5), ZN => n_138);
  g24027 : NR2XD0BWP7T port map(A1 => n_303, A2 => n_181, ZN => n_461);
  g24029 : NR2XD0BWP7T port map(A1 => n_424, A2 => n_181, ZN => n_220);
  g24000 : IND4D0BWP7T port map(A1 => ready, B1 => n_93, B2 => n_178, B3 => n_150, ZN => n_88);
  g24004 : INVD0BWP7T port map(I => n_433, ZN => n_86);
  g24008 : INVD0BWP7T port map(I => n_309, ZN => n_85);
  g24023 : ND4D0BWP7T port map(A1 => n_74, A2 => n_23, A3 => n_4, A4 => n_5, ZN => n_110);
  g23991 : NR2XD0BWP7T port map(A1 => n_78, A2 => n_96, ZN => n_95);
  g24015 : NR2XD0BWP7T port map(A1 => n_49, A2 => n_1589, ZN => n_92);
  g24021 : INVD1BWP7T port map(I => n_84, ZN => n_306);
  g24032 : INVD1BWP7T port map(I => n_83, ZN => n_274);
  g24006 : INVD1BWP7T port map(I => n_82, ZN => n_368);
  g24033 : INVD0BWP7T port map(I => n_356, ZN => n_81);
  g24051 : INVD0BWP7T port map(I => n_303, ZN => n_80);
  g24007 : INVD0BWP7T port map(I => n_326, ZN => n_79);
  g24035 : INVD1BWP7T port map(I => n_424, ZN => n_180);
  g23993 : NR2XD0BWP7T port map(A1 => n_78, A2 => counter(1), ZN => n_91);
  g24036 : INVD0BWP7T port map(I => n_149, ZN => n_134);
  g24034 : INVD1BWP7T port map(I => n_77, ZN => n_388);
  g24049 : INVD1BWP7T port map(I => n_76, ZN => n_340);
  g24048 : INVD1BWP7T port map(I => n_75, ZN => n_280);
  g24050 : INVD1BWP7T port map(I => n_182, ZN => n_405);
  g24031 : INR2D1BWP7T port map(A1 => n_71, B1 => n_72, ZN => n_84);
  g24042 : INR2D1BWP7T port map(A1 => n_74, B1 => n_1589, ZN => n_83);
  g24016 : NR2XD0BWP7T port map(A1 => n_72, A2 => n_1589, ZN => n_82);
  g24026 : ND3D0BWP7T port map(A1 => n_71, A2 => n_53, A3 => counter(4), ZN => n_97);
  g24039 : ND2D1BWP7T port map(A1 => n_70, A2 => n_69, ZN => n_151);
  g24038 : IND2D0BWP7T port map(A1 => n_119, B1 => counter(4), ZN => n_117);
  g24040 : ND2D1BWP7T port map(A1 => n_29, A2 => state(0), ZN => n_148);
  g24020 : INVD1BWP7T port map(I => n_68, ZN => n_284);
  g24041 : ND2D0BWP7T port map(A1 => n_155, A2 => sqi_finished, ZN => n_161);
  g24018 : ND2D1BWP7T port map(A1 => n_67, A2 => n_58, ZN => n_309);
  g24017 : ND2D1BWP7T port map(A1 => n_67, A2 => n_71, ZN => n_326);
  g24044 : NR2D0BWP7T port map(A1 => n_63, A2 => n_1589, ZN => n_77);
  g24059 : INR2XD0BWP7T port map(A1 => n_59, B1 => n_63, ZN => n_76);
  g24055 : OA21D0BWP7T port map(A1 => n_62, A2 => n_2, B => ready, Z => n_105);
  g24058 : NR2D0BWP7T port map(A1 => n_63, A2 => n_52, ZN => n_75);
  g24060 : INR2XD0BWP7T port map(A1 => n_71, B1 => n_63, ZN => n_182);
  g24046 : INR2XD0BWP7T port map(A1 => n_61, B1 => n_104, ZN => n_149);
  g24009 : INVD1BWP7T port map(I => n_60, ZN => n_335);
  g24014 : ND2D1BWP7T port map(A1 => n_67, A2 => n_59, ZN => n_433);
  g24043 : ND2D1BWP7T port map(A1 => n_74, A2 => n_59, ZN => n_356);
  g24045 : ND2D1BWP7T port map(A1 => n_74, A2 => n_58, ZN => n_424);
  g24061 : ND2D1BWP7T port map(A1 => n_74, A2 => n_71, ZN => n_303);
  g24053 : AOI21D0BWP7T port map(A1 => n_181, A2 => n_93, B => n_99, ZN => n_56);
  g24074 : INVD0BWP7T port map(I => n_54, ZN => n_55);
  g24022 : ND3D0BWP7T port map(A1 => n_58, A2 => n_53, A3 => counter(4), ZN => n_78);
  g24030 : INR2XD0BWP7T port map(A1 => n_59, B1 => n_72, ZN => n_68);
  g24078 : INVD0BWP7T port map(I => n_155, ZN => n_94);
  g24019 : NR2XD0BWP7T port map(A1 => n_72, A2 => n_52, ZN => n_60);
  g24047 : INVD0BWP7T port map(I => n_67, ZN => n_49);
  g24037 : ND2D1BWP7T port map(A1 => n_150, A2 => sqi_finished, ZN => n_46);
  g24011 : IND2D1BWP7T port map(A1 => n_44, B1 => mode, ZN => n_45);
  g24025 : NR4D0BWP7T port map(A1 => n_17, A2 => counter(6), A3 => counter(5), A4 => counter(7), ZN => n_98);
  g24075 : INVD0BWP7T port map(I => n_100, ZN => n_36);
  g24062 : AN2D0BWP7T port map(A1 => n_34, A2 => n_93, Z => n_35);
  g24063 : NR2D0BWP7T port map(A1 => n_34, A2 => state(0), ZN => n_104);
  g24064 : IND2D0BWP7T port map(A1 => n_114, B1 => counter(3), ZN => n_119);
  g24065 : IND2D1BWP7T port map(A1 => n_33, B1 => n_13, ZN => n_63);
  g24057 : NR3D0BWP7T port map(A1 => n_33, A2 => n_32, A3 => counter(5), ZN => n_67);
  g24066 : NR2XD0BWP7T port map(A1 => n_27, A2 => counter(1), ZN => n_74);
  g24067 : ND2D1BWP7T port map(A1 => n_31, A2 => sqi_data_in(6), ZN => n_432);
  g24068 : ND2D1BWP7T port map(A1 => n_31, A2 => sqi_data_in(7), ZN => n_423);
  g24072 : ND2D1BWP7T port map(A1 => n_31, A2 => sqi_data_in(4), ZN => n_427);
  g24073 : ND2D1BWP7T port map(A1 => n_31, A2 => sqi_data_in(1), ZN => n_413);
  g24069 : ND2D1BWP7T port map(A1 => n_31, A2 => sqi_data_in(2), ZN => n_409);
  g24070 : ND2D1BWP7T port map(A1 => n_31, A2 => sqi_data_in(0), ZN => n_419);
  g24071 : ND2D1BWP7T port map(A1 => n_31, A2 => sqi_data_in(5), ZN => n_436);
  g24077 : INVD0BWP7T port map(I => n_150, ZN => n_30);
  g24079 : OAI21D0BWP7T port map(A1 => n_0, A2 => state(1), B => n_34, ZN => n_29);
  g24082 : ND2D1BWP7T port map(A1 => n_101, A2 => n_99, ZN => n_54);
  g24080 : IND3D1BWP7T port map(A1 => n_27, B1 => n_122, B2 => n_12, ZN => n_70);
  g24084 : ND2D4BWP7T port map(A1 => n_102, A2 => n_141, ZN => ready);
  g24087 : AN2D1BWP7T port map(A1 => n_23, A2 => sqi_finished, Z => n_71);
  g24090 : ND2D0BWP7T port map(A1 => n_181, A2 => n_184, ZN => n_155);
  g24091 : ND2D1BWP7T port map(A1 => n_31, A2 => sqi_data_in(3), ZN => n_402);
  g24092 : INVD0BWP7T port map(I => n_102, ZN => n_62);
  g24094 : INVD0BWP7T port map(I => n_178, ZN => n_69);
  g24054 : OAI211D1BWP7T port map(A1 => reset, A2 => n_141, B => ce, C => rw, ZN => n_44);
  g24081 : IND3D1BWP7T port map(A1 => state(2), B1 => state(3), B2 => n_18, ZN => n_61);
  g24083 : NR4D0BWP7T port map(A1 => n_1, A2 => x(4), A3 => x(0), A4 => x(1), ZN => n_100);
  g24076 : INVD1BWP7T port map(I => n_52, ZN => n_58);
  g24056 : ND4D0BWP7T port map(A1 => n_14, A2 => n_96, A3 => n_22, A4 => counter(3), ZN => n_72);
  g24107 : INVD0BWP7T port map(I => n_191, ZN => n_21);
  g24161 : INVD1BWP7T port map(I => reset, ZN => n_26);
  g24093 : INVD0BWP7T port map(I => n_181, ZN => n_65);
  g24146 : INVD1BWP7T port map(I => reset, ZN => n_2);
  g24168 : INVD1BWP7T port map(I => reset, ZN => n_25);
  g24086 : NR3D0BWP7T port map(A1 => n_9, A2 => counter(0), A3 => n_99, ZN => n_59);
  g24089 : IND3D1BWP7T port map(A1 => state(3), B1 => state(2), B2 => n_18, ZN => n_150);
  g24109 : AOI21D0BWP7T port map(A1 => n_32, A2 => n_16, B => n_15, ZN => n_17);
  g24101 : ND2D1BWP7T port map(A1 => n_14, A2 => n_13, ZN => n_27);
  g24095 : INR2D1BWP7T port map(A1 => n_13, B1 => counter(7), ZN => n_53);
  g24088 : ND3D0BWP7T port map(A1 => n_12, A2 => counter(0), A3 => sqi_finished, ZN => n_52);
  g24108 : INVD1BWP7T port map(I => n_184, ZN => n_31);
  g24106 : OR2D1BWP7T port map(A1 => n_7, A2 => state(0), Z => n_178);
  g24105 : ND2D1BWP7T port map(A1 => n_18, A2 => n_8, ZN => n_181);
  g24112 : ND2D1BWP7T port map(A1 => n_14, A2 => counter(1), ZN => n_33);
  g24102 : AN2D0BWP7T port map(A1 => n_12, A2 => n_144, Z => n_23);
  g24114 : IND2D0BWP7T port map(A1 => n_122, B1 => counter(2), ZN => n_114);
  g24113 : ND2D1BWP7T port map(A1 => n_8, A2 => state(1), ZN => n_34);
  g24104 : IND2D1BWP7T port map(A1 => n_6, B1 => state(0), ZN => n_102);
  g24116 : ND2D1BWP7T port map(A1 => n_8, A2 => state(0), ZN => n_93);
  g24115 : IND2D1BWP7T port map(A1 => n_7, B1 => state(0), ZN => n_101);
  g24117 : NR2D1BWP7T port map(A1 => n_6, A2 => state(0), ZN => n_191);
  g24110 : NR4D0BWP7T port map(A1 => y(2), A2 => y(0), A3 => y(4), A4 => y(6), ZN => n_5);
  g24111 : NR4D0BWP7T port map(A1 => y(3), A2 => y(1), A3 => y(5), A4 => y(7), ZN => n_4);
  g24120 : ND2D1BWP7T port map(A1 => n_137, A2 => counter(2), ZN => n_9);
  g24118 : IND3D1BWP7T port map(A1 => state(1), B1 => state(2), B2 => state(0), ZN => n_184);
  g24126 : CKND2D1BWP7T port map(A1 => state(1), A2 => state(2), ZN => n_7);
  g24123 : NR2XD0BWP7T port map(A1 => counter(4), A2 => counter(7), ZN => n_14);
  g24128 : NR2XD0BWP7T port map(A1 => counter(3), A2 => counter(5), ZN => n_13);
  g24122 : NR2XD0BWP7T port map(A1 => counter(2), A2 => counter(6), ZN => n_12);
  g24130 : CKND2D1BWP7T port map(A1 => counter(0), A2 => counter(1), ZN => n_122);
  g24125 : OR2D1BWP7T port map(A1 => x(2), A2 => x(3), Z => n_1);
  g24127 : CKND2D1BWP7T port map(A1 => state(1), A2 => state(3), ZN => n_6);
  g24129 : NR2D1BWP7T port map(A1 => state(2), A2 => state(3), ZN => n_8);
  g24121 : NR2D1BWP7T port map(A1 => state(1), A2 => state(0), ZN => n_18);
  g24124 : CKND2D1BWP7T port map(A1 => state(2), A2 => state(3), ZN => n_141);
  g24132 : INVD1BWP7T port map(I => sqi_finished, ZN => n_99);
  g2 : ND2D1BWP7T port map(A1 => n_65, A2 => sqi_finished, ZN => n_493);
  drc_bufs24402 : INVD4BWP7T port map(I => n_496, ZN => framebuffer_buf(0));
  drc_bufs24408 : INVD4BWP7T port map(I => n_502, ZN => framebuffer_buf(157));
  drc_bufs24414 : INVD4BWP7T port map(I => n_508, ZN => framebuffer_buf(156));
  drc_bufs24420 : INVD4BWP7T port map(I => n_514, ZN => framebuffer_buf(7));
  drc_bufs24426 : INVD4BWP7T port map(I => n_520, ZN => framebuffer_buf(154));
  drc_bufs24432 : INVD4BWP7T port map(I => n_526, ZN => framebuffer_buf(153));
  drc_bufs24438 : INVD4BWP7T port map(I => n_532, ZN => framebuffer_buf(152));
  drc_bufs24444 : INVD4BWP7T port map(I => n_538, ZN => framebuffer_buf(8));
  drc_bufs24450 : INVD4BWP7T port map(I => n_544, ZN => framebuffer_buf(150));
  drc_bufs24456 : INVD4BWP7T port map(I => n_550, ZN => framebuffer_buf(149));
  drc_bufs24462 : INVD4BWP7T port map(I => n_556, ZN => framebuffer_buf(148));
  drc_bufs24468 : INVD4BWP7T port map(I => n_562, ZN => framebuffer_buf(147));
  drc_bufs24474 : INVD4BWP7T port map(I => n_568, ZN => framebuffer_buf(146));
  drc_bufs24480 : INVD4BWP7T port map(I => n_574, ZN => framebuffer_buf(145));
  drc_bufs24486 : INVD4BWP7T port map(I => n_580, ZN => framebuffer_buf(144));
  drc_bufs24492 : INVD4BWP7T port map(I => n_586, ZN => framebuffer_buf(9));
  drc_bufs24498 : INVD4BWP7T port map(I => n_592, ZN => framebuffer_buf(142));
  drc_bufs24504 : INVD4BWP7T port map(I => n_598, ZN => framebuffer_buf(141));
  drc_bufs24510 : INVD4BWP7T port map(I => n_604, ZN => framebuffer_buf(140));
  drc_bufs24516 : INVD4BWP7T port map(I => n_610, ZN => framebuffer_buf(39));
  drc_bufs24522 : INVD4BWP7T port map(I => n_616, ZN => framebuffer_buf(138));
  drc_bufs24528 : INVD4BWP7T port map(I => n_622, ZN => framebuffer_buf(40));
  drc_bufs24534 : INVD4BWP7T port map(I => n_628, ZN => framebuffer_buf(136));
  drc_bufs24540 : INVD4BWP7T port map(I => n_634, ZN => framebuffer_buf(103));
  drc_bufs24546 : INVD4BWP7T port map(I => n_640, ZN => framebuffer_buf(134));
  drc_bufs24552 : INVD4BWP7T port map(I => n_646, ZN => framebuffer_buf(133));
  drc_bufs24558 : INVD4BWP7T port map(I => n_652, ZN => framebuffer_buf(132));
  drc_bufs24564 : INVD4BWP7T port map(I => n_658, ZN => framebuffer_buf(131));
  drc_bufs24570 : INVD4BWP7T port map(I => n_664, ZN => framebuffer_buf(130));
  drc_bufs24576 : INVD4BWP7T port map(I => n_670, ZN => framebuffer_buf(129));
  drc_bufs24582 : INVD4BWP7T port map(I => n_676, ZN => framebuffer_buf(128));
  drc_bufs24588 : INVD4BWP7T port map(I => n_682, ZN => framebuffer_buf(104));
  drc_bufs24594 : INVD4BWP7T port map(I => n_688, ZN => framebuffer_buf(126));
  drc_bufs24600 : INVD4BWP7T port map(I => n_694, ZN => framebuffer_buf(125));
  drc_bufs24606 : INVD4BWP7T port map(I => n_700, ZN => framebuffer_buf(124));
  drc_bufs24612 : INVD4BWP7T port map(I => n_706, ZN => framebuffer_buf(105));
  drc_bufs24618 : INVD4BWP7T port map(I => n_712, ZN => framebuffer_buf(122));
  drc_bufs24624 : INVD4BWP7T port map(I => n_718, ZN => framebuffer_buf(121));
  drc_bufs24630 : INVD4BWP7T port map(I => n_724, ZN => framebuffer_buf(120));
  drc_bufs24636 : INVD4BWP7T port map(I => n_730, ZN => framebuffer_buf(106));
  drc_bufs24642 : INVD4BWP7T port map(I => n_736, ZN => framebuffer_buf(118));
  drc_bufs24648 : INVD4BWP7T port map(I => n_742, ZN => framebuffer_buf(117));
  drc_bufs24654 : INVD4BWP7T port map(I => n_748, ZN => framebuffer_buf(116));
  drc_bufs24660 : INVD4BWP7T port map(I => n_754, ZN => framebuffer_buf(41));
  drc_bufs24666 : INVD4BWP7T port map(I => n_760, ZN => framebuffer_buf(114));
  drc_bufs24672 : INVD4BWP7T port map(I => n_766, ZN => framebuffer_buf(113));
  drc_bufs24678 : INVD4BWP7T port map(I => n_772, ZN => framebuffer_buf(112));
  drc_bufs24684 : INVD4BWP7T port map(I => n_778, ZN => framebuffer_buf(107));
  drc_bufs24690 : INVD4BWP7T port map(I => n_784, ZN => framebuffer_buf(108));
  drc_bufs24696 : INVD4BWP7T port map(I => n_790, ZN => framebuffer_buf(42));
  drc_bufs24702 : INVD4BWP7T port map(I => n_796, ZN => framebuffer_buf(109));
  drc_bufs24708 : INVD4BWP7T port map(I => n_802, ZN => framebuffer_buf(110));
  drc_bufs24714 : INVD4BWP7T port map(I => n_808, ZN => framebuffer_buf(10));
  drc_bufs24720 : INVD4BWP7T port map(I => n_814, ZN => framebuffer_buf(43));
  drc_bufs24726 : INVD4BWP7T port map(I => n_820, ZN => framebuffer_buf(111));
  drc_bufs24732 : INVD4BWP7T port map(I => n_826, ZN => framebuffer_buf(44));
  drc_bufs24738 : INVD4BWP7T port map(I => n_832, ZN => framebuffer_buf(102));
  drc_bufs24744 : INVD4BWP7T port map(I => n_838, ZN => framebuffer_buf(101));
  drc_bufs24750 : INVD4BWP7T port map(I => n_844, ZN => framebuffer_buf(100));
  drc_bufs24756 : INVD4BWP7T port map(I => n_850, ZN => framebuffer_buf(99));
  drc_bufs24762 : INVD4BWP7T port map(I => n_856, ZN => framebuffer_buf(98));
  drc_bufs24768 : INVD4BWP7T port map(I => n_862, ZN => framebuffer_buf(97));
  drc_bufs24774 : INVD4BWP7T port map(I => n_868, ZN => framebuffer_buf(96));
  drc_bufs24780 : INVD4BWP7T port map(I => n_874, ZN => framebuffer_buf(45));
  drc_bufs24786 : INVD4BWP7T port map(I => n_880, ZN => framebuffer_buf(94));
  drc_bufs24792 : INVD4BWP7T port map(I => n_886, ZN => framebuffer_buf(93));
  drc_bufs24798 : INVD4BWP7T port map(I => n_892, ZN => framebuffer_buf(92));
  drc_bufs24804 : INVD4BWP7T port map(I => n_898, ZN => framebuffer_buf(115));
  drc_bufs24810 : INVD4BWP7T port map(I => n_904, ZN => framebuffer_buf(90));
  drc_bufs24816 : INVD4BWP7T port map(I => n_910, ZN => framebuffer_buf(89));
  drc_bufs24822 : INVD4BWP7T port map(I => n_916, ZN => framebuffer_buf(88));
  drc_bufs24828 : INVD4BWP7T port map(I => n_922, ZN => framebuffer_buf(46));
  drc_bufs24834 : INVD4BWP7T port map(I => n_928, ZN => framebuffer_buf(86));
  drc_bufs24840 : INVD4BWP7T port map(I => n_934, ZN => framebuffer_buf(85));
  drc_bufs24846 : INVD4BWP7T port map(I => n_940, ZN => framebuffer_buf(84));
  drc_bufs24852 : INVD4BWP7T port map(I => n_946, ZN => framebuffer_buf(11));
  drc_bufs24858 : INVD4BWP7T port map(I => n_952, ZN => framebuffer_buf(82));
  drc_bufs24864 : INVD4BWP7T port map(I => n_958, ZN => framebuffer_buf(12));
  drc_bufs24870 : INVD4BWP7T port map(I => n_964, ZN => framebuffer_buf(80));
  drc_bufs24876 : INVD4BWP7T port map(I => n_970, ZN => framebuffer_buf(47));
  drc_bufs24882 : INVD4BWP7T port map(I => n_976, ZN => framebuffer_buf(78));
  drc_bufs24888 : INVD4BWP7T port map(I => n_982, ZN => framebuffer_buf(77));
  drc_bufs24894 : INVD4BWP7T port map(I => n_988, ZN => framebuffer_buf(76));
  drc_bufs24900 : INVD4BWP7T port map(I => n_994, ZN => framebuffer_buf(119));
  drc_bufs24906 : INVD4BWP7T port map(I => n_1000, ZN => framebuffer_buf(74));
  drc_bufs24912 : INVD4BWP7T port map(I => n_1006, ZN => framebuffer_buf(48));
  drc_bufs24918 : INVD4BWP7T port map(I => n_1012, ZN => framebuffer_buf(72));
  drc_bufs24924 : INVD4BWP7T port map(I => n_1018, ZN => framebuffer_buf(49));
  drc_bufs24930 : INVD4BWP7T port map(I => n_1024, ZN => framebuffer_buf(70));
  drc_bufs24936 : INVD4BWP7T port map(I => n_1030, ZN => framebuffer_buf(69));
  drc_bufs24942 : INVD4BWP7T port map(I => n_1036, ZN => framebuffer_buf(68));
  drc_bufs24948 : INVD4BWP7T port map(I => n_1042, ZN => framebuffer_buf(123));
  drc_bufs24954 : INVD4BWP7T port map(I => n_1048, ZN => framebuffer_buf(66));
  drc_bufs24960 : INVD4BWP7T port map(I => n_1054, ZN => framebuffer_buf(155));
  drc_bufs24966 : INVD4BWP7T port map(I => n_1060, ZN => framebuffer_buf(64));
  drc_bufs24972 : INVD4BWP7T port map(I => n_1066, ZN => framebuffer_buf(151));
  drc_bufs24978 : INVD4BWP7T port map(I => n_1072, ZN => framebuffer_buf(62));
  drc_bufs24984 : INVD4BWP7T port map(I => n_1078, ZN => framebuffer_buf(61));
  drc_bufs24990 : INVD4BWP7T port map(I => n_1084, ZN => framebuffer_buf(60));
  drc_bufs24996 : INVD4BWP7T port map(I => n_1090, ZN => framebuffer_buf(143));
  drc_bufs25002 : INVD4BWP7T port map(I => n_1096, ZN => framebuffer_buf(58));
  drc_bufs25008 : INVD4BWP7T port map(I => n_1102, ZN => framebuffer_buf(139));
  drc_bufs25014 : INVD4BWP7T port map(I => n_1108, ZN => framebuffer_buf(137));
  drc_bufs25020 : INVD4BWP7T port map(I => n_1114, ZN => framebuffer_buf(135));
  drc_bufs25026 : INVD4BWP7T port map(I => n_1120, ZN => framebuffer_buf(54));
  drc_bufs25032 : INVD4BWP7T port map(I => n_1126, ZN => framebuffer_buf(53));
  drc_bufs25038 : INVD4BWP7T port map(I => n_1132, ZN => framebuffer_buf(50));
  drc_bufs25044 : INVD4BWP7T port map(I => n_1138, ZN => framebuffer_buf(13));
  drc_bufs25050 : INVD4BWP7T port map(I => n_1144, ZN => framebuffer_buf(51));
  drc_bufs25056 : INVD4BWP7T port map(I => n_1150, ZN => framebuffer_buf(127));
  drc_bufs25062 : INVD4BWP7T port map(I => n_1156, ZN => framebuffer_buf(52));
  drc_bufs25068 : INVD4BWP7T port map(I => n_1162, ZN => framebuffer_buf(14));
  drc_bufs25074 : INVD4BWP7T port map(I => n_1168, ZN => framebuffer_buf(15));
  drc_bufs25080 : INVD4BWP7T port map(I => n_1174, ZN => framebuffer_buf(16));
  drc_bufs25086 : INVD4BWP7T port map(I => n_1180, ZN => framebuffer_buf(55));
  drc_bufs25092 : INVD4BWP7T port map(I => n_1186, ZN => framebuffer_buf(56));
  drc_bufs25098 : INVD4BWP7T port map(I => n_1192, ZN => framebuffer_buf(57));
  drc_bufs25104 : INVD4BWP7T port map(I => n_1198, ZN => framebuffer_buf(17));
  drc_bufs25110 : INVD4BWP7T port map(I => n_1204, ZN => framebuffer_buf(59));
  drc_bufs25116 : INVD4BWP7T port map(I => n_1210, ZN => framebuffer_buf(18));
  drc_bufs25122 : INVD4BWP7T port map(I => n_1216, ZN => framebuffer_buf(38));
  drc_bufs25128 : INVD4BWP7T port map(I => n_1222, ZN => framebuffer_buf(37));
  drc_bufs25134 : INVD4BWP7T port map(I => n_1228, ZN => framebuffer_buf(36));
  drc_bufs25140 : INVD4BWP7T port map(I => n_1234, ZN => framebuffer_buf(95));
  drc_bufs25146 : INVD4BWP7T port map(I => n_1240, ZN => framebuffer_buf(34));
  drc_bufs25152 : INVD4BWP7T port map(I => n_1246, ZN => framebuffer_buf(91));
  drc_bufs25158 : INVD4BWP7T port map(I => n_1252, ZN => framebuffer_buf(32));
  drc_bufs25164 : INVD4BWP7T port map(I => n_1258, ZN => framebuffer_buf(87));
  drc_bufs25170 : INVD4BWP7T port map(I => n_1264, ZN => framebuffer_buf(30));
  drc_bufs25176 : INVD4BWP7T port map(I => n_1270, ZN => framebuffer_buf(83));
  drc_bufs25182 : INVD4BWP7T port map(I => n_1276, ZN => framebuffer_buf(81));
  drc_bufs25188 : INVD4BWP7T port map(I => n_1282, ZN => framebuffer_buf(79));
  drc_bufs25194 : INVD4BWP7T port map(I => n_1288, ZN => framebuffer_buf(26));
  drc_bufs25200 : INVD4BWP7T port map(I => n_1294, ZN => framebuffer_buf(75));
  drc_bufs25206 : INVD4BWP7T port map(I => n_1300, ZN => framebuffer_buf(73));
  drc_bufs25212 : INVD4BWP7T port map(I => n_1306, ZN => framebuffer_buf(71));
  drc_bufs25218 : INVD4BWP7T port map(I => n_1312, ZN => framebuffer_buf(22));
  drc_bufs25224 : INVD4BWP7T port map(I => n_1318, ZN => framebuffer_buf(67));
  drc_bufs25230 : INVD4BWP7T port map(I => n_1324, ZN => framebuffer_buf(19));
  drc_bufs25236 : INVD4BWP7T port map(I => n_1330, ZN => framebuffer_buf(20));
  drc_bufs25242 : INVD4BWP7T port map(I => n_1336, ZN => framebuffer_buf(63));
  drc_bufs25248 : INVD4BWP7T port map(I => n_1342, ZN => framebuffer_buf(65));
  drc_bufs25254 : INVD4BWP7T port map(I => n_1348, ZN => framebuffer_buf(21));
  drc_bufs25260 : INVD4BWP7T port map(I => n_1354, ZN => framebuffer_buf(1));
  drc_bufs25266 : INVD4BWP7T port map(I => n_1360, ZN => framebuffer_buf(2));
  drc_bufs25272 : INVD4BWP7T port map(I => n_1366, ZN => framebuffer_buf(23));
  drc_bufs25278 : INVD4BWP7T port map(I => n_1372, ZN => framebuffer_buf(24));
  drc_bufs25284 : INVD4BWP7T port map(I => n_1378, ZN => framebuffer_buf(25));
  drc_bufs25290 : INVD4BWP7T port map(I => n_1384, ZN => framebuffer_buf(27));
  drc_bufs25296 : INVD4BWP7T port map(I => n_1390, ZN => framebuffer_buf(28));
  drc_bufs25302 : INVD4BWP7T port map(I => n_1396, ZN => framebuffer_buf(29));
  drc_bufs25308 : INVD4BWP7T port map(I => n_1402, ZN => framebuffer_buf(3));
  drc_bufs25314 : INVD4BWP7T port map(I => n_1408, ZN => framebuffer_buf(6));
  drc_bufs25320 : INVD4BWP7T port map(I => n_1414, ZN => framebuffer_buf(35));
  drc_bufs25326 : INVD4BWP7T port map(I => n_1422, ZN => framebuffer_buf(4));
  drc_bufs25332 : INVD4BWP7T port map(I => n_1428, ZN => framebuffer_buf(31));
  drc_bufs25338 : INVD4BWP7T port map(I => n_1434, ZN => framebuffer_buf(33));
  drc_bufs25344 : INVD4BWP7T port map(I => n_1440, ZN => framebuffer_buf(5));
  drc_bufs25350 : INVD4BWP7T port map(I => n_1446, ZN => calc_buf_out(23));
  drc_bufs25356 : INVD4BWP7T port map(I => n_1452, ZN => calc_buf_out(6));
  drc_bufs25362 : INVD4BWP7T port map(I => n_1458, ZN => calc_buf_out(9));
  drc_bufs25368 : INVD4BWP7T port map(I => n_1464, ZN => calc_buf_out(21));
  drc_bufs25374 : INVD4BWP7T port map(I => n_1470, ZN => calc_buf_out(1));
  drc_bufs25380 : INVD4BWP7T port map(I => n_1476, ZN => calc_buf_out(20));
  drc_bufs25386 : INVD4BWP7T port map(I => n_1482, ZN => calc_buf_out(12));
  drc_bufs25392 : INVD4BWP7T port map(I => n_1488, ZN => calc_buf_out(5));
  drc_bufs25398 : INVD4BWP7T port map(I => n_1494, ZN => calc_buf_out(15));
  drc_bufs25404 : INVD4BWP7T port map(I => n_1500, ZN => calc_buf_out(17));
  drc_bufs25410 : INVD4BWP7T port map(I => n_1506, ZN => calc_buf_out(16));
  drc_bufs25416 : INVD4BWP7T port map(I => n_1512, ZN => calc_buf_out(4));
  drc_bufs25422 : INVD4BWP7T port map(I => n_1518, ZN => calc_buf_out(10));
  drc_bufs25428 : INVD4BWP7T port map(I => n_1524, ZN => calc_buf_out(22));
  drc_bufs25434 : INVD4BWP7T port map(I => n_1530, ZN => calc_buf_out(8));
  drc_bufs25440 : INVD4BWP7T port map(I => n_1536, ZN => calc_buf_out(18));
  drc_bufs25446 : INVD4BWP7T port map(I => n_1542, ZN => calc_buf_out(0));
  drc_bufs25452 : INVD4BWP7T port map(I => n_1548, ZN => calc_buf_out(14));
  drc_bufs25458 : INVD4BWP7T port map(I => n_1554, ZN => calc_buf_out(2));
  drc_bufs25464 : INVD4BWP7T port map(I => n_1560, ZN => calc_buf_out(7));
  drc_bufs25470 : INVD4BWP7T port map(I => n_1566, ZN => calc_buf_out(19));
  drc_bufs25476 : INVD4BWP7T port map(I => n_1572, ZN => calc_buf_out(13));
  drc_bufs25482 : INVD4BWP7T port map(I => n_1578, ZN => calc_buf_out(11));
  drc_bufs25488 : INVD4BWP7T port map(I => n_1584, ZN => calc_buf_out(3));
  state_reg_3 : DFD1BWP7T port map(CP => clk, D => n_152, Q => state(3), QN => n_0);
  counter_reg_3 : DFKCND1BWP7T port map(CP => clk, CN => n_2, D => new_counter(3), Q => counter(3), QN => n_32);
  counter_reg_0 : DFKCND1BWP7T port map(CP => clk, CN => n_2, D => new_counter(0), Q => counter(0), QN => n_144);
  counter_reg_1 : DFKCND1BWP7T port map(CP => clk, CN => n_2, D => new_counter(1), Q => counter(1), QN => n_96);
  counter_reg_5 : DFKCND1BWP7T port map(CP => clk, CN => n_2, D => new_counter(5), Q => counter(5), QN => n_22);
  counter_reg_2 : DFKCND1BWP7T port map(CP => clk, CN => n_2, D => new_counter(2), Q => counter(2), QN => n_16);
  counter_reg_4 : DFKCND1BWP7T port map(CP => clk, CN => n_2, D => new_counter(4), Q => counter(4), QN => n_15);
  counter_reg_6 : DFKCND1BWP7T port map(CP => clk, CN => n_2, D => new_counter(6), Q => counter(6), QN => n_137);
  framebuffer_buf_reg_0 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_311, Q => framebuffer_buf_0_2333, QN => n_496);
  framebuffer_buf_reg_157 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_354, Q => framebuffer_buf_157_2490, QN => n_502);
  framebuffer_buf_reg_156 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_358, Q => framebuffer_buf_156_2489, QN => n_508);
  framebuffer_buf_reg_7 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_238, Q => framebuffer_buf_7_2340, QN => n_514);
  framebuffer_buf_reg_154 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_361, Q => framebuffer_buf_154_2487, QN => n_520);
  framebuffer_buf_reg_153 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_364, Q => framebuffer_buf_153_2486, QN => n_526);
  framebuffer_buf_reg_152 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_366, Q => framebuffer_buf_152_2485, QN => n_532);
  framebuffer_buf_reg_8 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_237, Q => framebuffer_buf_8_2341, QN => n_538);
  framebuffer_buf_reg_150 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_373, Q => framebuffer_buf_150_2483, QN => n_544);
  framebuffer_buf_reg_149 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_374, Q => framebuffer_buf_149_2482, QN => n_550);
  framebuffer_buf_reg_148 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_376, Q => framebuffer_buf_148_2481, QN => n_556);
  framebuffer_buf_reg_147 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_377, Q => framebuffer_buf_147_2480, QN => n_562);
  framebuffer_buf_reg_146 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_378, Q => framebuffer_buf_146_2479, QN => n_568);
  framebuffer_buf_reg_145 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_382, Q => framebuffer_buf_145_2478, QN => n_574);
  framebuffer_buf_reg_144 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_384, Q => framebuffer_buf_144_2477, QN => n_580);
  framebuffer_buf_reg_9 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_235, Q => framebuffer_buf_9_2342, QN => n_586);
  framebuffer_buf_reg_142 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_352, Q => framebuffer_buf_142_2475, QN => n_592);
  framebuffer_buf_reg_141 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_398, Q => framebuffer_buf_141_2474, QN => n_598);
  framebuffer_buf_reg_140 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_400, Q => framebuffer_buf_140_2473, QN => n_604);
  framebuffer_buf_reg_39 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_344, Q => framebuffer_buf_39_2372, QN => n_610);
  framebuffer_buf_reg_138 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_410, Q => framebuffer_buf_138_2471, QN => n_616);
  framebuffer_buf_reg_40 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_270, Q => framebuffer_buf_40_2373, QN => n_622);
  framebuffer_buf_reg_136 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_421, Q => framebuffer_buf_136_2469, QN => n_628);
  framebuffer_buf_reg_103 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_240, Q => framebuffer_buf_103_2436, QN => n_634);
  framebuffer_buf_reg_134 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_365, Q => framebuffer_buf_134_2467, QN => n_640);
  framebuffer_buf_reg_133 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_437, Q => framebuffer_buf_133_2466, QN => n_646);
  framebuffer_buf_reg_132 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_429, Q => framebuffer_buf_132_2465, QN => n_652);
  framebuffer_buf_reg_131 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_224, Q => framebuffer_buf_131_2464, QN => n_658);
  framebuffer_buf_reg_130 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_228, Q => framebuffer_buf_130_2463, QN => n_664);
  framebuffer_buf_reg_129 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_230, Q => framebuffer_buf_129_2462, QN => n_670);
  framebuffer_buf_reg_128 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_236, Q => framebuffer_buf_128_2461, QN => n_676);
  framebuffer_buf_reg_104 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_251, Q => framebuffer_buf_104_2437, QN => n_682);
  framebuffer_buf_reg_126 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_397, Q => framebuffer_buf_126_2459, QN => n_688);
  framebuffer_buf_reg_125 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_399, Q => framebuffer_buf_125_2458, QN => n_694);
  framebuffer_buf_reg_124 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_401, Q => framebuffer_buf_124_2457, QN => n_700);
  framebuffer_buf_reg_105 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_248, Q => framebuffer_buf_105_2438, QN => n_706);
  framebuffer_buf_reg_122 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_411, Q => framebuffer_buf_122_2455, QN => n_712);
  framebuffer_buf_reg_121 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_418, Q => framebuffer_buf_121_2454, QN => n_718);
  framebuffer_buf_reg_120 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_420, Q => framebuffer_buf_120_2453, QN => n_724);
  framebuffer_buf_reg_106 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_245, Q => framebuffer_buf_106_2439, QN => n_730);
  framebuffer_buf_reg_118 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_434, Q => framebuffer_buf_118_2451, QN => n_736);
  framebuffer_buf_reg_117 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_438, Q => framebuffer_buf_117_2450, QN => n_742);
  framebuffer_buf_reg_116 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_268, Q => framebuffer_buf_116_2449, QN => n_748);
  framebuffer_buf_reg_41 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_275, Q => framebuffer_buf_41_2374, QN => n_754);
  framebuffer_buf_reg_114 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_227, Q => framebuffer_buf_114_2447, QN => n_760);
  framebuffer_buf_reg_113 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_229, Q => framebuffer_buf_113_2446, QN => n_766);
  framebuffer_buf_reg_112 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_233, Q => framebuffer_buf_112_2445, QN => n_772);
  framebuffer_buf_reg_107 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_242, Q => framebuffer_buf_107_2440, QN => n_778);
  framebuffer_buf_reg_108 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_239, Q => framebuffer_buf_108_2441, QN => n_784);
  framebuffer_buf_reg_42 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_277, Q => framebuffer_buf_42_2375, QN => n_790);
  framebuffer_buf_reg_109 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_232, Q => framebuffer_buf_109_2442, QN => n_796);
  framebuffer_buf_reg_110 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_371, Q => framebuffer_buf_110_2443, QN => n_802);
  framebuffer_buf_reg_10 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_234, Q => framebuffer_buf_10_2343, QN => n_808);
  framebuffer_buf_reg_43 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_266, Q => framebuffer_buf_43_2376, QN => n_814);
  framebuffer_buf_reg_111 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_369, Q => framebuffer_buf_111_2444, QN => n_820);
  framebuffer_buf_reg_44 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_263, Q => framebuffer_buf_44_2377, QN => n_826);
  framebuffer_buf_reg_102 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_241, Q => framebuffer_buf_102_2435, QN => n_832);
  framebuffer_buf_reg_101 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_244, Q => framebuffer_buf_101_2434, QN => n_838);
  framebuffer_buf_reg_100 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_247, Q => framebuffer_buf_100_2433, QN => n_844);
  framebuffer_buf_reg_99 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_249, Q => framebuffer_buf_99_2432, QN => n_850);
  framebuffer_buf_reg_98 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_250, Q => framebuffer_buf_98_2431, QN => n_856);
  framebuffer_buf_reg_97 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_285, Q => framebuffer_buf_97_2430, QN => n_862);
  framebuffer_buf_reg_96 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_291, Q => framebuffer_buf_96_2429, QN => n_868);
  framebuffer_buf_reg_45 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_260, Q => framebuffer_buf_45_2378, QN => n_874);
  framebuffer_buf_reg_94 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_294, Q => framebuffer_buf_94_2427, QN => n_880);
  framebuffer_buf_reg_93 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_295, Q => framebuffer_buf_93_2426, QN => n_886);
  framebuffer_buf_reg_92 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_296, Q => framebuffer_buf_92_2425, QN => n_892);
  framebuffer_buf_reg_115 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_225, Q => framebuffer_buf_115_2448, QN => n_898);
  framebuffer_buf_reg_90 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_300, Q => framebuffer_buf_90_2423, QN => n_904);
  framebuffer_buf_reg_89 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_310, Q => framebuffer_buf_89_2422, QN => n_910);
  framebuffer_buf_reg_88 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_312, Q => framebuffer_buf_88_2421, QN => n_916);
  framebuffer_buf_reg_46 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_254, Q => framebuffer_buf_46_2379, QN => n_922);
  framebuffer_buf_reg_86 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_316, Q => framebuffer_buf_86_2419, QN => n_928);
  framebuffer_buf_reg_85 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_318, Q => framebuffer_buf_85_2418, QN => n_934);
  framebuffer_buf_reg_84 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_439, Q => framebuffer_buf_84_2417, QN => n_940);
  framebuffer_buf_reg_11 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_231, Q => framebuffer_buf_11_2344, QN => n_946);
  framebuffer_buf_reg_82 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_322, Q => framebuffer_buf_82_2415, QN => n_952);
  framebuffer_buf_reg_12 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_226, Q => framebuffer_buf_12_2345, QN => n_958);
  framebuffer_buf_reg_80 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_327, Q => framebuffer_buf_80_2413, QN => n_964);
  framebuffer_buf_reg_47 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_252, Q => framebuffer_buf_47_2380, QN => n_970);
  framebuffer_buf_reg_78 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_321, Q => framebuffer_buf_78_2411, QN => n_976);
  framebuffer_buf_reg_77 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_317, Q => framebuffer_buf_77_2410, QN => n_982);
  framebuffer_buf_reg_76 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_324, Q => framebuffer_buf_76_2409, QN => n_988);
  framebuffer_buf_reg_119 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_430, Q => framebuffer_buf_119_2452, QN => n_994);
  framebuffer_buf_reg_74 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_333, Q => framebuffer_buf_74_2407, QN => n_1000);
  framebuffer_buf_reg_48 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_343, Q => framebuffer_buf_48_2381, QN => n_1006);
  framebuffer_buf_reg_72 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_342, Q => framebuffer_buf_72_2405, QN => n_1012);
  framebuffer_buf_reg_49 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_341, Q => framebuffer_buf_49_2382, QN => n_1018);
  framebuffer_buf_reg_70 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_288, Q => framebuffer_buf_70_2403, QN => n_1024);
  framebuffer_buf_reg_69 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_290, Q => framebuffer_buf_69_2402, QN => n_1030);
  framebuffer_buf_reg_68 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_293, Q => framebuffer_buf_68_2401, QN => n_1036);
  framebuffer_buf_reg_123 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_407, Q => framebuffer_buf_123_2456, QN => n_1042);
  framebuffer_buf_reg_66 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_301, Q => framebuffer_buf_66_2399, QN => n_1048);
  framebuffer_buf_reg_155 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_360, Q => framebuffer_buf_155_2488, QN => n_1054);
  framebuffer_buf_reg_64 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_313, Q => framebuffer_buf_64_2397, QN => n_1060);
  framebuffer_buf_reg_151 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_372, Q => framebuffer_buf_151_2484, QN => n_1066);
  framebuffer_buf_reg_62 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_348, Q => framebuffer_buf_62_2395, QN => n_1072);
  framebuffer_buf_reg_61 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_375, Q => framebuffer_buf_61_2394, QN => n_1078);
  framebuffer_buf_reg_60 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_379, Q => framebuffer_buf_60_2393, QN => n_1084);
  framebuffer_buf_reg_143 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_350, Q => framebuffer_buf_143_2476, QN => n_1090);
  framebuffer_buf_reg_58 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_385, Q => framebuffer_buf_58_2391, QN => n_1096);
  framebuffer_buf_reg_139 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_403, Q => framebuffer_buf_139_2472, QN => n_1102);
  framebuffer_buf_reg_137 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_415, Q => framebuffer_buf_137_2470, QN => n_1108);
  framebuffer_buf_reg_135 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_359, Q => framebuffer_buf_135_2468, QN => n_1114);
  framebuffer_buf_reg_54 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_329, Q => framebuffer_buf_54_2387, QN => n_1120);
  framebuffer_buf_reg_53 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_331, Q => framebuffer_buf_53_2386, QN => n_1126);
  framebuffer_buf_reg_50 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_338, Q => framebuffer_buf_50_2383, QN => n_1132);
  framebuffer_buf_reg_13 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_319, Q => framebuffer_buf_13_2346, QN => n_1138);
  framebuffer_buf_reg_51 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_337, Q => framebuffer_buf_51_2384, QN => n_1144);
  framebuffer_buf_reg_127 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_394, Q => framebuffer_buf_127_2460, QN => n_1150);
  framebuffer_buf_reg_52 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_332, Q => framebuffer_buf_52_2385, QN => n_1156);
  framebuffer_buf_reg_14 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_435, Q => framebuffer_buf_14_2347, QN => n_1162);
  framebuffer_buf_reg_15 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_425, Q => framebuffer_buf_15_2348, QN => n_1168);
  framebuffer_buf_reg_16 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_408, Q => framebuffer_buf_16_2349, QN => n_1174);
  framebuffer_buf_reg_55 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_328, Q => framebuffer_buf_55_2388, QN => n_1180);
  framebuffer_buf_reg_56 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_395, Q => framebuffer_buf_56_2389, QN => n_1186);
  framebuffer_buf_reg_57 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_389, Q => framebuffer_buf_57_2390, QN => n_1192);
  framebuffer_buf_reg_17 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_406, Q => framebuffer_buf_17_2350, QN => n_1198);
  framebuffer_buf_reg_59 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_383, Q => framebuffer_buf_59_2392, QN => n_1204);
  framebuffer_buf_reg_18 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_396, Q => framebuffer_buf_18_2351, QN => n_1210);
  framebuffer_buf_reg_38 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_345, Q => framebuffer_buf_38_2371, QN => n_1216);
  framebuffer_buf_reg_37 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_347, Q => framebuffer_buf_37_2370, QN => n_1222);
  framebuffer_buf_reg_36 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_349, Q => framebuffer_buf_36_2369, QN => n_1228);
  framebuffer_buf_reg_95 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_292, Q => framebuffer_buf_95_2428, QN => n_1234);
  framebuffer_buf_reg_34 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_353, Q => framebuffer_buf_34_2367, QN => n_1240);
  framebuffer_buf_reg_91 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_299, Q => framebuffer_buf_91_2424, QN => n_1246);
  framebuffer_buf_reg_32 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_370, Q => framebuffer_buf_32_2365, QN => n_1252);
  framebuffer_buf_reg_87 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_314, Q => framebuffer_buf_87_2420, QN => n_1258);
  framebuffer_buf_reg_30 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_258, Q => framebuffer_buf_30_2363, QN => n_1264);
  framebuffer_buf_reg_83 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_320, Q => framebuffer_buf_83_2416, QN => n_1270);
  framebuffer_buf_reg_81 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_323, Q => framebuffer_buf_81_2414, QN => n_1276);
  framebuffer_buf_reg_79 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_315, Q => framebuffer_buf_79_2412, QN => n_1282);
  framebuffer_buf_reg_26 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_278, Q => framebuffer_buf_26_2359, QN => n_1288);
  framebuffer_buf_reg_75 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_330, Q => framebuffer_buf_75_2408, QN => n_1294);
  framebuffer_buf_reg_73 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_336, Q => framebuffer_buf_73_2406, QN => n_1300);
  framebuffer_buf_reg_71 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_286, Q => framebuffer_buf_71_2404, QN => n_1306);
  framebuffer_buf_reg_22 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_390, Q => framebuffer_buf_22_2355, QN => n_1312);
  framebuffer_buf_reg_67 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_297, Q => framebuffer_buf_67_2400, QN => n_1318);
  framebuffer_buf_reg_19 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_393, Q => framebuffer_buf_19_2352, QN => n_1324);
  framebuffer_buf_reg_20 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_392, Q => framebuffer_buf_20_2353, QN => n_1330);
  framebuffer_buf_reg_63 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_346, Q => framebuffer_buf_63_2396, QN => n_1336);
  framebuffer_buf_reg_65 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_307, Q => framebuffer_buf_65_2398, QN => n_1342);
  framebuffer_buf_reg_21 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_391, Q => framebuffer_buf_21_2354, QN => n_1348);
  framebuffer_buf_reg_1 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_304, Q => framebuffer_buf_1_2334, QN => n_1354);
  framebuffer_buf_reg_2 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_298, Q => framebuffer_buf_2_2335, QN => n_1360);
  framebuffer_buf_reg_23 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_386, Q => framebuffer_buf_23_2356, QN => n_1366);
  framebuffer_buf_reg_24 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_282, Q => framebuffer_buf_24_2357, QN => n_1372);
  framebuffer_buf_reg_25 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_281, Q => framebuffer_buf_25_2358, QN => n_1378);
  framebuffer_buf_reg_27 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_276, Q => framebuffer_buf_27_2360, QN => n_1384);
  framebuffer_buf_reg_28 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_272, Q => framebuffer_buf_28_2361, QN => n_1390);
  framebuffer_buf_reg_29 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_271, Q => framebuffer_buf_29_2362, QN => n_1396);
  framebuffer_buf_reg_3 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_289, Q => framebuffer_buf_3_2336, QN => n_1402);
  framebuffer_buf_reg_6 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_243, Q => framebuffer_buf_6_2339, QN => n_1408);
  framebuffer_buf_reg_35 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_351, Q => framebuffer_buf_35_2368, QN => n_1414);
  framebuffer_buf_reg_4 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_287, Q => framebuffer_buf_4_2337, QN => n_1422);
  framebuffer_buf_reg_31 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_256, Q => framebuffer_buf_31_2364, QN => n_1428);
  framebuffer_buf_reg_33 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_357, Q => framebuffer_buf_33_2366, QN => n_1434);
  framebuffer_buf_reg_5 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_246, Q => framebuffer_buf_5_2338, QN => n_1440);
  calc_buf_out_reg_23 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_218, Q => calc_buf_out_23_2332, QN => n_1446);
  calc_buf_out_reg_6 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_445, Q => calc_buf_out_6_2315, QN => n_1452);
  calc_buf_out_reg_9 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_223, Q => calc_buf_out_9_2318, QN => n_1458);
  calc_buf_out_reg_21 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_206, Q => calc_buf_out_21_2330, QN => n_1464);
  calc_buf_out_reg_1 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_444, Q => calc_buf_out_1_2310, QN => n_1470);
  calc_buf_out_reg_20 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_213, Q => calc_buf_out_20_2329, QN => n_1476);
  calc_buf_out_reg_12 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_215, Q => calc_buf_out_12_2321, QN => n_1482);
  calc_buf_out_reg_5 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_463, Q => calc_buf_out_5_2314, QN => n_1488);
  calc_buf_out_reg_15 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_214, Q => calc_buf_out_15_2324, QN => n_1494);
  calc_buf_out_reg_17 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_210, Q => calc_buf_out_17_2326, QN => n_1500);
  calc_buf_out_reg_16 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_207, Q => calc_buf_out_16_2325, QN => n_1506);
  calc_buf_out_reg_4 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_459, Q => calc_buf_out_4_2313, QN => n_1512);
  calc_buf_out_reg_10 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_216, Q => calc_buf_out_10_2319, QN => n_1518);
  calc_buf_out_reg_22 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_205, Q => calc_buf_out_22_2331, QN => n_1524);
  calc_buf_out_reg_8 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_204, Q => calc_buf_out_8_2317, QN => n_1530);
  calc_buf_out_reg_18 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_209, Q => calc_buf_out_18_2327, QN => n_1536);
  calc_buf_out_reg_0 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_443, Q => calc_buf_out_0_2309, QN => n_1542);
  calc_buf_out_reg_14 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_217, Q => calc_buf_out_14_2323, QN => n_1548);
  calc_buf_out_reg_2 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_462, Q => calc_buf_out_2_2311, QN => n_1554);
  calc_buf_out_reg_7 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_446, Q => calc_buf_out_7_2316, QN => n_1560);
  calc_buf_out_reg_19 : DFKCND0BWP7T port map(CP => clk, CN => n_2, D => n_208, Q => calc_buf_out_19_2328, QN => n_1566);
  calc_buf_out_reg_13 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_222, Q => calc_buf_out_13_2322, QN => n_1572);
  calc_buf_out_reg_11 : DFKCND0BWP7T port map(CP => clk, CN => n_26, D => n_219, Q => calc_buf_out_11_2320, QN => n_1578);
  calc_buf_out_reg_3 : DFKCND0BWP7T port map(CP => clk, CN => n_25, D => n_460, Q => calc_buf_out_3_2312, QN => n_1584);
  g25873 : IND4D0BWP7T port map(A1 => n_135, B1 => n_149, B2 => n_150, B3 => n_102, ZN => n_1588);
  g25874 : IND3D1BWP7T port map(A1 => n_9, B1 => counter(0), B2 => sqi_finished, ZN => n_1589);

end synthesised;
