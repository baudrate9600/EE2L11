configuration memory_behaviour_cfg of memory is
   for behaviour
   end for;
end memory_behaviour_cfg;
