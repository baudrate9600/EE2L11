library IEEE;
use IEEE.std_logic_1164.ALL;

entity test is
   port(test : in  std_logic);
end test;

