configuration tri_buffer_behaviour_cfg of tri_buffer is
   for behaviour
   end for;
end tri_buffer_behaviour_cfg;
