configuration memory_routed_cfg of memory is
   for routed
   end for;
end memory_routed_cfg;
