library IEEE;
use IEEE.std_logic_1164.ALL;

entity sram_test_tb is
end sram_test_tb;

