configuration address_alu_behaviour_cfg of address_alu is
   for behaviour
   end for;
end address_alu_behaviour_cfg;
