configuration shift_register_routed_cfg of shift_register is
   for routed
   end for;
end shift_register_routed_cfg;
