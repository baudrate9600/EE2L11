configuration sqi_controller_routed_cfg of sqi_controller is
   for routed
   end for;
end sqi_controller_routed_cfg;
