configuration line_buffer_behaviour_cfg of line_buffer is
   for behaviour
   end for;
end line_buffer_behaviour_cfg;
