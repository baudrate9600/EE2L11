configuration memory_tb_synthesised_behaviour_cfg of memory_tb is
   for behaviour
      for all: memory use configuration work.memory_synthesised_cfg;
      end for;
   end for;
end memory_tb_synthesised_behaviour_cfg;
