configuration sqi_routed_cfg of sqi is
   for routed
   end for;
end sqi_routed_cfg;
