configuration sqi_behaviour_cfg of sqi is
   for behaviour
   end for;
end sqi_behaviour_cfg;
