library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.all; 
architecture behaviour of abs_address is
begin
		process(reg) is begin

	  end process; 
end behaviour;

