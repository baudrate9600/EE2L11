configuration shift_register_synthesised_cfg of shift_register is
   for synthesised
   end for;
end shift_register_synthesised_cfg;
