configuration sram_interface_synthesised_cfg of sram_interface is
   for synthesised
   end for;
end sram_interface_synthesised_cfg;
