configuration counter16_synthesised_cfg of counter16 is
   for synthesised
   end for;
end counter16_synthesised_cfg;
