LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
ARCHITECTURE behaviour OF sqi IS
 	SIGNAL count_reset: std_logic;
	SIGNAL count_en   : std_logic;
	SIGNAL count_load : std_logic;
	SIGNAL count_in   : std_logic_vector(3 DOWNTO 0);
	SIGNAL count_out  : std_logic_vector(3 DOWNTO 0);
 

	SIGNAL data_wire  : std_logic_vector(7 DOWNTO 0);
	SIGNAL data_read  : std_logic_vector(7 DOWNTO 0); 
	SIGNAL data_read_in: std_logic_vector (7 DOWNTO 0); 

	SIGNAL load_reg   : std_logic;
	SIGNAL shift_reg  : std_logic;
	SIGNAL shift_in   : std_logic_vector(3 DOWNTO 0);
	SIGNAL shift_out  : std_logic_vector(3 DOWNTO 0);
  SIGNAL shift_reset : std_logic; 

	SIGNAL mux_select : std_logic_vector(2 DOWNTO 0); 

	SIGNAL spi_wire   : std_logic;
 
	--All the components
	COMPONENT counter16 IS
		PORT 
		(
			clk       : IN std_logic;
			reset     : IN std_logic;
			load      : IN std_logic;
			enable    : IN std_logic;
			count_in  : IN std_logic_vector(3 DOWNTO 0);
			count_out : OUT std_logic_vector(3 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT shift_register IS
		PORT 
		(
			clk       : IN std_logic;
			reset     : IN std_logic;
			load      : IN std_logic;
			shift     : IN std_logic;
			data_in   : IN std_logic_vector(7 DOWNTO 0);
			data_out  : OUT std_logic_vector(7 DOWNTO 0);
			shift_in  : IN std_logic_vector(3 DOWNTO 0);
			shift_out : OUT std_logic_vector(3 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT sqi_controller IS
		PORT 
		(
			clk      : IN std_logic;
			reset    : IN std_logic;
			en       : IN std_logic;
			RW       : IN std_logic;
			high_z 		: OUT std_logic; 
			new_data : OUT std_logic; 
			single			: IN std_logic; 
			data_in  : IN std_logic_vector(7 DOWNTO 0);
			shift_data_in    : in std_logic_vector(7 downto 0);
			data_read: OUT std_logic_vector(7 downto 0);
			data_out : OUT std_logic_vector(7 DOWNTO 0);
			address  : IN std_logic_vector(14 DOWNTO 0);
			--counter interface
			count_reset: OUT std_logic;
			count_en   : OUT std_logic;
			count_load : OUT std_logic;
			count_in   : IN std_logic_vector(3 DOWNTO 0);
			count_out  : OUT std_logic_vector(3 DOWNTO 0);
			--shift register interface
			reg_shift : OUT std_logic;
			reg_load  : OUT std_logic;
			done      : OUT std_logic;
			shift_in  : IN std_logic_vector(3 DOWNTO 0);
			shift_reset : OUT std_logic;
			--SQI wires
			sck  : OUT std_logic;
			cs   : OUT std_logic;
			MOSI : OUT std_logic_vector (3 DOWNTO 0)
		);
	END COMPONENT;

BEGIN
	u0 : counter16
	PORT MAP(clk, count_reset, count_load, count_en, count_in, count_out);
	u1 : shift_register
	PORT MAP(clk, shift_reset, load_reg, shift_reg, data_wire, data_read_in, MISO, shift_out);
	u2 : sqi_controller
	PORT MAP
	(clk,reset,en,RW,high_z,new_data,single,data_in,data_read_in, data_out,data_wire,address,count_reset,count_en,count_load,count_out,count_in, 
		shift_reg,load_reg,done,shift_out,shift_reset,SCK,CS,MOSI );

 
 
 
END behaviour;

