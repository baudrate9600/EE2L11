library IEEE;
use IEEE.std_logic_1164.ALL;

entity address_alu_tb is
end address_alu_tb;

