configuration sqi_tb_behaviour_cfg2 of sqi_tb is
   for behaviour
      for all: sqi use configuration work.sqi_routed_cfg;
      end for;
   end for;
end sqi_tb_behaviour_cfg2;
