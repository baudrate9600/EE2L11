
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture routed of memory is

  component DEL01BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD5BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL1BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD4BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD12BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD6BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component INVD2BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component DFKCNQD1BWP7T
    port(CN, CP, D : in std_logic; Q : out std_logic);
  end component;

  component LHQD1BWP7T
    port(D, E : in std_logic; Q : out std_logic);
  end component;

  component AO32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component OAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD5BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component NR3D1BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component LHD1BWP7T
    port(D, E : in std_logic; Q, QN : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OR4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI211XD0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component IND3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component LNQD1BWP7T
    port(D, EN : in std_logic; Q : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OA211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component NR4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CN, CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component DFKCND0BWP7T
    port(CN, CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  signal FE_PHN188_framebuffer_buf_10_2298, FE_PHN187_framebuffer_buf_104_2392, FE_PHN186_framebuffer_buf_14_2302, FE_PHN185_framebuffer_buf_153_2441, FE_PHN184_framebuffer_buf_150_2438 : std_logic;
  signal FE_PHN183_framebuffer_buf_66_2354, FE_PHN182_framebuffer_buf_92_2380, FE_PHN181_framebuffer_buf_39_2327, FE_PHN180_framebuffer_buf_105_2393, FE_PHN179_framebuffer_buf_123_2411 : std_logic;
  signal FE_PHN178_framebuffer_buf_118_2406, FE_PHN177_framebuffer_buf_151_2439, FE_PHN176_calc_buf_out_20_2284, FE_PHN175_framebuffer_buf_109_2397, FE_PHN174_framebuffer_buf_20_2308 : std_logic;
  signal FE_PHN173_framebuffer_buf_39_2327, FE_PHN172_framebuffer_buf_134_2422, FE_PHN171_framebuffer_buf_44_2332, FE_PHN170_framebuffer_buf_131_2419, FE_PHN169_calc_buf_out_20_2284 : std_logic;
  signal FE_PHN168_framebuffer_buf_56_2344, FE_PHN167_framebuffer_buf_130_2418, FE_PHN166_framebuffer_buf_1_2289, FE_PHN165_framebuffer_buf_50_2338, FE_PHN164_framebuffer_buf_129_2417 : std_logic;
  signal FE_PHN163_framebuffer_buf_93_2381, FE_PHN162_framebuffer_buf_151_2439, FE_PHN161_framebuffer_buf_136_2424, FE_PHN160_framebuffer_buf_10_2298, FE_PHN159_framebuffer_buf_150_2438 : std_logic;
  signal FE_PHN158_framebuffer_buf_117_2405, FE_PHN157_framebuffer_buf_104_2392, FE_PHN156_framebuffer_buf_143_2431, FE_PHN155_framebuffer_buf_138_2426, FE_PHN154_framebuffer_buf_105_2393 : std_logic;
  signal FE_PHN153_framebuffer_buf_108_2396, FE_PHN152_framebuffer_buf_43_2331, FE_PHN151_framebuffer_buf_75_2363, FE_PHN150_calc_buf_out_21_2285, FE_PHN149_framebuffer_buf_118_2406 : std_logic;
  signal FE_PHN148_framebuffer_buf_78_2366, FE_PHN147_framebuffer_buf_32_2320, FE_PHN146_framebuffer_buf_107_2395, FE_PHN145_framebuffer_buf_84_2372, FE_PHN144_framebuffer_buf_23_2311 : std_logic;
  signal FE_PHN143_framebuffer_buf_14_2302, FE_PHN142_framebuffer_buf_62_2350, FE_PHN141_calc_buf_out_19_2283, FE_PHN140_framebuffer_buf_42_2330, FE_PHN139_framebuffer_buf_153_2441 : std_logic;
  signal FE_PHN138_framebuffer_buf_60_2348, FE_PHN137_framebuffer_buf_80_2368, FE_PHN136_framebuffer_buf_71_2359, FE_PHN135_framebuffer_buf_47_2335, FE_PHN134_framebuffer_buf_99_2387 : std_logic;
  signal FE_PHN133_framebuffer_buf_21_2309, FE_PHN132_framebuffer_buf_28_2316, FE_PHN131_framebuffer_buf_16_2304, FE_PHN130_framebuffer_buf_92_2380, FE_PHN129_framebuffer_buf_26_2314 : std_logic;
  signal FE_PHN128_framebuffer_buf_29_2317, FE_PHN127_framebuffer_buf_123_2411, FE_PHN126_framebuffer_buf_8_2296, FE_PHN125_framebuffer_buf_114_2402, FE_PHN124_framebuffer_buf_73_2361 : std_logic;
  signal FE_PHN123_framebuffer_buf_35_2323, FE_PHN122_framebuffer_buf_12_2300, FE_PHN121_framebuffer_buf_3_2291, FE_PHN120_framebuffer_buf_31_2319, FE_PHN119_framebuffer_buf_66_2354 : std_logic;
  signal FE_PHN118_framebuffer_buf_154_2442, FE_PHN117_framebuffer_buf_102_2390, FE_PHN116_framebuffer_buf_55_2343, FE_PHN115_framebuffer_buf_27_2315, FE_PHN114_framebuffer_buf_85_2373 : std_logic;
  signal FE_PHN113_framebuffer_buf_37_2325, FE_PHN112_framebuffer_buf_25_2313, FE_PHN111_framebuffer_buf_113_2401, FE_PHN110_calc_buf_out_15_2279, FE_PHN109_framebuffer_buf_46_2334 : std_logic;
  signal FE_PHN108_framebuffer_buf_126_2414, FE_PHN107_framebuffer_buf_135_2423, FE_PHN106_framebuffer_buf_59_2347, FE_PHN105_framebuffer_buf_145_2433, FE_PHN104_framebuffer_buf_36_2324 : std_logic;
  signal FE_PHN103_framebuffer_buf_34_2322, FE_PHN102_framebuffer_buf_81_2369, FE_PHN101_framebuffer_buf_5_2293, FE_PHN100_framebuffer_buf_86_2374, FE_PHN99_framebuffer_buf_137_2425 : std_logic;
  signal FE_PHN98_framebuffer_buf_98_2386, FE_PHN97_framebuffer_buf_156_2444, FE_PHN96_framebuffer_buf_124_2412, FE_PHN95_framebuffer_buf_38_2326, FE_PHN94_framebuffer_buf_140_2428 : std_logic;
  signal FE_PHN93_calc_buf_out_12_2276, FE_PHN92_framebuffer_buf_7_2295, FE_PHN91_framebuffer_buf_132_2420, FE_PHN90_framebuffer_buf_45_2333, FE_PHN89_framebuffer_buf_88_2376 : std_logic;
  signal FE_PHN88_framebuffer_buf_139_2427, FE_PHN87_framebuffer_buf_142_2430, FE_PHN86_framebuffer_buf_54_2342, FE_PHN85_framebuffer_buf_48_2336, FE_PHN84_framebuffer_buf_70_2358 : std_logic;
  signal FE_PHN83_framebuffer_buf_33_2321, FE_PHN82_framebuffer_buf_24_2312, FE_PHN81_framebuffer_buf_76_2364, FE_PHN80_framebuffer_buf_146_2434, FE_PHN79_framebuffer_buf_91_2379 : std_logic;
  signal FE_PHN78_framebuffer_buf_63_2351, FE_PHN77_framebuffer_buf_17_2305, FE_PHN76_framebuffer_buf_30_2318, FE_PHN75_framebuffer_buf_120_2408, FE_PHN74_framebuffer_buf_116_2404 : std_logic;
  signal FE_PHN73_framebuffer_buf_52_2340, FE_PHN72_framebuffer_buf_87_2375, FE_PHN71_framebuffer_buf_111_2399, FE_PHN70_framebuffer_buf_100_2388, FE_PHN69_framebuffer_buf_2_2290 : std_logic;
  signal FE_PHN68_framebuffer_buf_9_2297, FE_PHN67_framebuffer_buf_6_2294, FE_PHN66_framebuffer_buf_41_2329, FE_PHN65_framebuffer_buf_125_2413, FE_PHN64_framebuffer_buf_64_2352 : std_logic;
  signal FE_PHN63_framebuffer_buf_95_2383, FE_PHN62_framebuffer_buf_94_2382, FE_PHN61_calc_buf_out_23_2287, FE_PHN60_framebuffer_buf_0_2288, FE_PHN59_framebuffer_buf_112_2400 : std_logic;
  signal FE_PHN58_framebuffer_buf_51_2339, FE_PHN57_framebuffer_buf_58_2346, FE_PHN56_framebuffer_buf_103_2391, FE_PHN55_framebuffer_buf_101_2389, FE_PHN54_framebuffer_buf_96_2384 : std_logic;
  signal FE_PHN53_framebuffer_buf_69_2357, FE_PHN52_framebuffer_buf_110_2398, FE_PHN51_framebuffer_buf_128_2416, FE_PHN50_framebuffer_buf_4_2292, FE_PHN49_framebuffer_buf_141_2429 : std_logic;
  signal FE_PHN48_framebuffer_buf_72_2360, FE_PHN47_framebuffer_buf_106_2394, FE_PHN46_framebuffer_buf_97_2385, FE_PHN45_framebuffer_buf_122_2410, FE_PHN44_framebuffer_buf_157_2445 : std_logic;
  signal FE_PHN43_framebuffer_buf_53_2341, FE_PHN42_framebuffer_buf_19_2307, FE_PHN41_calc_buf_out_16_2280, FE_PHN40_framebuffer_buf_61_2349, FE_PHN39_calc_buf_out_10_2274 : std_logic;
  signal FE_PHN38_framebuffer_buf_144_2432, FE_PHN37_calc_buf_out_13_2277, FE_PHN36_framebuffer_buf_119_2407, FE_PHN35_calc_buf_out_9_2273, FE_PHN34_framebuffer_buf_68_2356 : std_logic;
  signal FE_PHN33_framebuffer_buf_11_2299, FE_PHN32_calc_buf_out_14_2278, FE_PHN31_framebuffer_buf_89_2377, FE_PHN30_framebuffer_buf_18_2306, FE_PHN29_framebuffer_buf_121_2409 : std_logic;
  signal FE_PHN28_calc_buf_out_22_2286, FE_PHN27_framebuffer_buf_127_2415, FE_PHN26_calc_buf_out_18_2282, FE_PHN25_calc_buf_out_11_2275, FE_PHN24_framebuffer_buf_155_2443 : std_logic;
  signal FE_PHN23_calc_buf_out_17_2281, FE_PHN22_calc_buf_out_8_2272, FE_PHN21_framebuffer_buf_149_2437, FE_PHN20_framebuffer_buf_79_2367, FE_PHN19_framebuffer_buf_15_2303 : std_logic;
  signal FE_PHN18_framebuffer_buf_22_2310, FE_PHN17_framebuffer_buf_74_2362, FE_PHN16_framebuffer_buf_65_2353, FE_PHN15_framebuffer_buf_77_2365, FE_PHN14_framebuffer_buf_13_2301 : std_logic;
  signal FE_PHN13_framebuffer_buf_148_2436, FE_PHN12_framebuffer_buf_67_2355, FE_PHN11_framebuffer_buf_57_2345, FE_PHN10_framebuffer_buf_83_2371, FE_PHN9_framebuffer_buf_90_2378 : std_logic;
  signal FE_PHN8_framebuffer_buf_49_2337, FE_PHN7_framebuffer_buf_152_2440, FE_PHN6_framebuffer_buf_133_2421, FE_PHN5_framebuffer_buf_82_2370, FE_PHN4_framebuffer_buf_115_2403 : std_logic;
  signal FE_PHN3_framebuffer_buf_40_2328, FE_PHN2_framebuffer_buf_147_2435, FE_OFN1_FE_DBTN0_reset, FE_OFN0_FE_DBTN0_reset, CTS_14 : std_logic;
  signal CTS_13, CTS_12, FE_DBTN0_reset : std_logic;
  signal new_counter : std_logic_vector(7 downto 0);
  signal counter : std_logic_vector(7 downto 0);
  signal new_calc_buf_out : std_logic_vector(23 downto 0);
  signal state : std_logic_vector(3 downto 0);
  signal row_buf : std_logic_vector(5 downto 0);
  signal new_row_buf : std_logic_vector(5 downto 0);
  signal UNCONNECTED, UNCONNECTED0, UNCONNECTED1, UNCONNECTED2, UNCONNECTED3 : std_logic;
  signal UNCONNECTED4, UNCONNECTED5, UNCONNECTED6, calc_buf_out_0_2264, calc_buf_out_1_2265 : std_logic;
  signal calc_buf_out_2_2266, calc_buf_out_3_2267, calc_buf_out_4_2268, calc_buf_out_5_2269, calc_buf_out_6_2270 : std_logic;
  signal calc_buf_out_7_2271, calc_buf_out_8_2272, calc_buf_out_9_2273, calc_buf_out_10_2274, calc_buf_out_11_2275 : std_logic;
  signal calc_buf_out_12_2276, calc_buf_out_13_2277, calc_buf_out_14_2278, calc_buf_out_15_2279, calc_buf_out_16_2280 : std_logic;
  signal calc_buf_out_17_2281, calc_buf_out_18_2282, calc_buf_out_19_2283, calc_buf_out_20_2284, calc_buf_out_21_2285 : std_logic;
  signal calc_buf_out_22_2286, calc_buf_out_23_2287, framebuffer_buf_0_2288, framebuffer_buf_1_2289, framebuffer_buf_2_2290 : std_logic;
  signal framebuffer_buf_3_2291, framebuffer_buf_4_2292, framebuffer_buf_5_2293, framebuffer_buf_6_2294, framebuffer_buf_7_2295 : std_logic;
  signal framebuffer_buf_8_2296, framebuffer_buf_9_2297, framebuffer_buf_10_2298, framebuffer_buf_11_2299, framebuffer_buf_12_2300 : std_logic;
  signal framebuffer_buf_13_2301, framebuffer_buf_14_2302, framebuffer_buf_15_2303, framebuffer_buf_16_2304, framebuffer_buf_17_2305 : std_logic;
  signal framebuffer_buf_18_2306, framebuffer_buf_19_2307, framebuffer_buf_20_2308, framebuffer_buf_21_2309, framebuffer_buf_22_2310 : std_logic;
  signal framebuffer_buf_23_2311, framebuffer_buf_24_2312, framebuffer_buf_25_2313, framebuffer_buf_26_2314, framebuffer_buf_27_2315 : std_logic;
  signal framebuffer_buf_28_2316, framebuffer_buf_29_2317, framebuffer_buf_30_2318, framebuffer_buf_31_2319, framebuffer_buf_32_2320 : std_logic;
  signal framebuffer_buf_33_2321, framebuffer_buf_34_2322, framebuffer_buf_35_2323, framebuffer_buf_36_2324, framebuffer_buf_37_2325 : std_logic;
  signal framebuffer_buf_38_2326, framebuffer_buf_39_2327, framebuffer_buf_40_2328, framebuffer_buf_41_2329, framebuffer_buf_42_2330 : std_logic;
  signal framebuffer_buf_43_2331, framebuffer_buf_44_2332, framebuffer_buf_45_2333, framebuffer_buf_46_2334, framebuffer_buf_47_2335 : std_logic;
  signal framebuffer_buf_48_2336, framebuffer_buf_49_2337, framebuffer_buf_50_2338, framebuffer_buf_51_2339, framebuffer_buf_52_2340 : std_logic;
  signal framebuffer_buf_53_2341, framebuffer_buf_54_2342, framebuffer_buf_55_2343, framebuffer_buf_56_2344, framebuffer_buf_57_2345 : std_logic;
  signal framebuffer_buf_58_2346, framebuffer_buf_59_2347, framebuffer_buf_60_2348, framebuffer_buf_61_2349, framebuffer_buf_62_2350 : std_logic;
  signal framebuffer_buf_63_2351, framebuffer_buf_64_2352, framebuffer_buf_65_2353, framebuffer_buf_66_2354, framebuffer_buf_67_2355 : std_logic;
  signal framebuffer_buf_68_2356, framebuffer_buf_69_2357, framebuffer_buf_70_2358, framebuffer_buf_71_2359, framebuffer_buf_72_2360 : std_logic;
  signal framebuffer_buf_73_2361, framebuffer_buf_74_2362, framebuffer_buf_75_2363, framebuffer_buf_76_2364, framebuffer_buf_77_2365 : std_logic;
  signal framebuffer_buf_78_2366, framebuffer_buf_79_2367, framebuffer_buf_80_2368, framebuffer_buf_81_2369, framebuffer_buf_82_2370 : std_logic;
  signal framebuffer_buf_83_2371, framebuffer_buf_84_2372, framebuffer_buf_85_2373, framebuffer_buf_86_2374, framebuffer_buf_87_2375 : std_logic;
  signal framebuffer_buf_88_2376, framebuffer_buf_89_2377, framebuffer_buf_90_2378, framebuffer_buf_91_2379, framebuffer_buf_92_2380 : std_logic;
  signal framebuffer_buf_93_2381, framebuffer_buf_94_2382, framebuffer_buf_95_2383, framebuffer_buf_96_2384, framebuffer_buf_97_2385 : std_logic;
  signal framebuffer_buf_98_2386, framebuffer_buf_99_2387, framebuffer_buf_100_2388, framebuffer_buf_101_2389, framebuffer_buf_102_2390 : std_logic;
  signal framebuffer_buf_103_2391, framebuffer_buf_104_2392, framebuffer_buf_105_2393, framebuffer_buf_106_2394, framebuffer_buf_107_2395 : std_logic;
  signal framebuffer_buf_108_2396, framebuffer_buf_109_2397, framebuffer_buf_110_2398, framebuffer_buf_111_2399, framebuffer_buf_112_2400 : std_logic;
  signal framebuffer_buf_113_2401, framebuffer_buf_114_2402, framebuffer_buf_115_2403, framebuffer_buf_116_2404, framebuffer_buf_117_2405 : std_logic;
  signal framebuffer_buf_118_2406, framebuffer_buf_119_2407, framebuffer_buf_120_2408, framebuffer_buf_121_2409, framebuffer_buf_122_2410 : std_logic;
  signal framebuffer_buf_123_2411, framebuffer_buf_124_2412, framebuffer_buf_125_2413, framebuffer_buf_126_2414, framebuffer_buf_127_2415 : std_logic;
  signal framebuffer_buf_128_2416, framebuffer_buf_129_2417, framebuffer_buf_130_2418, framebuffer_buf_131_2419, framebuffer_buf_132_2420 : std_logic;
  signal framebuffer_buf_133_2421, framebuffer_buf_134_2422, framebuffer_buf_135_2423, framebuffer_buf_136_2424, framebuffer_buf_137_2425 : std_logic;
  signal framebuffer_buf_138_2426, framebuffer_buf_139_2427, framebuffer_buf_140_2428, framebuffer_buf_141_2429, framebuffer_buf_142_2430 : std_logic;
  signal framebuffer_buf_143_2431, framebuffer_buf_144_2432, framebuffer_buf_145_2433, framebuffer_buf_146_2434, framebuffer_buf_147_2435 : std_logic;
  signal framebuffer_buf_148_2436, framebuffer_buf_149_2437, framebuffer_buf_150_2438, framebuffer_buf_151_2439, framebuffer_buf_152_2440 : std_logic;
  signal framebuffer_buf_153_2441, framebuffer_buf_154_2442, framebuffer_buf_155_2443, framebuffer_buf_156_2444, framebuffer_buf_157_2445 : std_logic;
  signal n_0, n_2, n_3, n_4, n_5 : std_logic;
  signal n_6, n_7, n_8, n_9, n_10 : std_logic;
  signal n_11, n_12, n_13, n_14, n_15 : std_logic;
  signal n_16, n_17, n_18, n_19, n_20 : std_logic;
  signal n_21, n_22, n_23, n_24, n_25 : std_logic;
  signal n_26, n_27, n_29, n_30, n_31 : std_logic;
  signal n_32, n_33, n_34, n_35, n_36 : std_logic;
  signal n_37, n_38, n_39, n_40, n_41 : std_logic;
  signal n_42, n_43, n_44, n_45, n_46 : std_logic;
  signal n_47, n_48, n_49, n_50, n_51 : std_logic;
  signal n_52, n_54, n_55, n_56, n_57 : std_logic;
  signal n_58, n_59, n_61, n_62, n_63 : std_logic;
  signal n_64, n_65, n_66, n_67, n_68 : std_logic;
  signal n_69, n_70, n_71, n_72, n_73 : std_logic;
  signal n_74, n_75, n_76, n_77, n_78 : std_logic;
  signal n_79, n_80, n_81, n_82, n_83 : std_logic;
  signal n_85, n_86, n_87, n_88, n_89 : std_logic;
  signal n_90, n_91, n_92, n_93, n_94 : std_logic;
  signal n_95, n_96, n_97, n_98, n_99 : std_logic;
  signal n_100, n_101, n_102, n_103, n_104 : std_logic;
  signal n_105, n_106, n_107, n_108, n_109 : std_logic;
  signal n_110, n_111, n_112, n_113, n_114 : std_logic;
  signal n_115, n_116, n_117, n_118, n_119 : std_logic;
  signal n_120, n_121, n_122, n_123, n_124 : std_logic;
  signal n_126, n_127, n_128, n_129, n_135 : std_logic;
  signal n_136, n_139, n_140, n_141, n_142 : std_logic;
  signal n_143, n_144, n_145, n_146, n_147 : std_logic;
  signal n_148, n_149, n_150, n_151, n_152 : std_logic;
  signal n_153, n_154, n_155, n_156, n_157 : std_logic;
  signal n_158, n_159, n_160, n_161, n_162 : std_logic;
  signal n_163, n_164, n_165, n_166, n_167 : std_logic;
  signal n_168, n_169, n_170, n_171, n_172 : std_logic;
  signal n_173, n_174, n_175, n_176, n_177 : std_logic;
  signal n_178, n_179, n_180, n_181, n_182 : std_logic;
  signal n_183, n_184, n_185, n_186, n_187 : std_logic;
  signal n_188, n_189, n_190, n_191, n_192 : std_logic;
  signal n_193, n_194, n_195, n_196, n_197 : std_logic;
  signal n_198, n_199, n_200, n_201, n_202 : std_logic;
  signal n_203, n_204, n_205, n_206, n_207 : std_logic;
  signal n_208, n_209, n_210, n_211, n_212 : std_logic;
  signal n_213, n_214, n_215, n_216, n_217 : std_logic;
  signal n_218, n_219, n_220, n_221, n_222 : std_logic;
  signal n_223, n_224, n_225, n_226, n_227 : std_logic;
  signal n_228, n_229, n_230, n_231, n_232 : std_logic;
  signal n_233, n_234, n_235, n_236, n_237 : std_logic;
  signal n_238, n_239, n_240, n_241, n_242 : std_logic;
  signal n_243, n_244, n_245, n_246, n_247 : std_logic;
  signal n_248, n_249, n_250, n_251, n_252 : std_logic;
  signal n_253, n_254, n_255, n_256, n_257 : std_logic;
  signal n_258, n_259, n_260, n_261, n_262 : std_logic;
  signal n_263, n_264, n_265, n_266, n_267 : std_logic;
  signal n_268, n_269, n_270, n_271, n_272 : std_logic;
  signal n_273, n_274, n_275, n_276, n_277 : std_logic;
  signal n_278, n_279, n_280, n_281, n_282 : std_logic;
  signal n_283, n_284, n_285, n_286, n_287 : std_logic;
  signal n_288, n_289, n_290, n_291, n_292 : std_logic;
  signal n_293, n_294, n_295, n_296, n_297 : std_logic;
  signal n_298, n_299, n_300, n_301, n_302 : std_logic;
  signal n_303, n_305, n_306, n_307, n_308 : std_logic;
  signal n_309, n_310, n_311, n_312, n_313 : std_logic;
  signal n_314, n_315, n_316, n_317, n_318 : std_logic;
  signal n_319, n_320, n_321, n_322, n_323 : std_logic;
  signal n_324, n_325, n_326, n_327, n_328 : std_logic;
  signal n_329, n_330, n_331, n_332, n_333 : std_logic;
  signal n_334, n_335, n_336, n_337, n_338 : std_logic;
  signal n_339, n_340, n_341, n_342, n_343 : std_logic;
  signal n_344, n_345, n_346, n_347, n_348 : std_logic;
  signal n_349, n_350, n_351, n_352, n_353 : std_logic;
  signal n_354, n_355, n_356, n_357, n_358 : std_logic;
  signal n_359, n_360, n_361, n_362, n_363 : std_logic;
  signal n_364, n_365, n_366, n_368, n_369 : std_logic;
  signal n_370, n_371, n_372, n_373, n_374 : std_logic;
  signal n_375, n_376, n_377, n_378, n_379 : std_logic;
  signal n_380, n_381, n_382, n_383, n_384 : std_logic;
  signal n_385, n_386, n_387, n_388, n_389 : std_logic;
  signal n_390, n_391, n_392, n_393, n_394 : std_logic;
  signal n_395, n_396, n_397, n_400, n_401 : std_logic;
  signal n_402, n_403, n_404, n_405, n_406 : std_logic;
  signal n_407, n_430, n_436, n_442, n_448 : std_logic;
  signal n_454, n_460, n_466, n_472, n_478 : std_logic;
  signal n_484, n_490, n_496, n_502, n_508 : std_logic;
  signal n_514, n_520, n_526, n_532, n_538 : std_logic;
  signal n_544, n_550, n_556, n_562, n_568 : std_logic;
  signal n_574, n_580, n_586, n_592, n_598 : std_logic;
  signal n_604, n_610, n_616, n_622, n_628 : std_logic;
  signal n_634, n_640, n_646, n_652, n_658 : std_logic;
  signal n_664, n_670, n_676, n_682, n_688 : std_logic;
  signal n_694, n_700, n_706, n_712, n_718 : std_logic;
  signal n_724, n_730, n_736, n_742, n_748 : std_logic;
  signal n_754, n_760, n_766, n_772, n_778 : std_logic;
  signal n_784, n_790, n_796, n_802, n_808 : std_logic;
  signal n_814, n_820, n_826, n_832, n_838 : std_logic;
  signal n_844, n_850, n_856, n_862, n_868 : std_logic;
  signal n_874, n_880, n_886, n_892, n_898 : std_logic;
  signal n_904, n_910, n_916, n_922, n_928 : std_logic;
  signal n_934, n_940, n_946, n_952, n_958 : std_logic;
  signal n_964, n_970, n_976, n_982, n_988 : std_logic;
  signal n_994, n_1000, n_1006, n_1012, n_1018 : std_logic;
  signal n_1024, n_1030, n_1036, n_1042, n_1048 : std_logic;
  signal n_1054, n_1060, n_1066, n_1072, n_1078 : std_logic;
  signal n_1084, n_1090, n_1096, n_1102, n_1108 : std_logic;
  signal n_1114, n_1120, n_1126, n_1132, n_1138 : std_logic;
  signal n_1144, n_1150, n_1156, n_1162, n_1168 : std_logic;
  signal n_1174, n_1180, n_1186, n_1192, n_1198 : std_logic;
  signal n_1204, n_1210, n_1216, n_1222, n_1228 : std_logic;
  signal n_1234, n_1240, n_1246, n_1252, n_1258 : std_logic;
  signal n_1264, n_1270, n_1276, n_1282, n_1288 : std_logic;
  signal n_1294, n_1300, n_1306, n_1312, n_1318 : std_logic;
  signal n_1324, n_1330, n_1336, n_1342, n_1348 : std_logic;
  signal n_1354, n_1362, n_1368, n_1374, n_1380 : std_logic;
  signal n_1386, n_1392, n_1398, n_1404, n_1410 : std_logic;
  signal n_1416, n_1422, n_1428, n_1434, n_1440 : std_logic;
  signal n_1446, n_1452, n_1458, n_1464, n_1470 : std_logic;
  signal n_1476, n_1482, n_1488, n_1494, n_1500 : std_logic;
  signal n_1506, n_1512, n_1518, n_1522, n_1523 : std_logic;

begin

  FE_PHC188_framebuffer_buf_10_2298 : DEL01BWP7T port map(I => FE_PHN160_framebuffer_buf_10_2298, Z => FE_PHN188_framebuffer_buf_10_2298);
  FE_PHC187_framebuffer_buf_104_2392 : DEL01BWP7T port map(I => FE_PHN187_framebuffer_buf_104_2392, Z => framebuffer_buf_104_2392);
  FE_PHC186_framebuffer_buf_14_2302 : DEL01BWP7T port map(I => FE_PHN186_framebuffer_buf_14_2302, Z => framebuffer_buf_14_2302);
  FE_PHC185_framebuffer_buf_153_2441 : DEL01BWP7T port map(I => FE_PHN139_framebuffer_buf_153_2441, Z => FE_PHN185_framebuffer_buf_153_2441);
  FE_PHC184_framebuffer_buf_150_2438 : DEL01BWP7T port map(I => FE_PHN184_framebuffer_buf_150_2438, Z => FE_PHN159_framebuffer_buf_150_2438);
  FE_PHC183_framebuffer_buf_66_2354 : DEL01BWP7T port map(I => FE_PHN119_framebuffer_buf_66_2354, Z => FE_PHN183_framebuffer_buf_66_2354);
  FE_PHC182_framebuffer_buf_92_2380 : DEL01BWP7T port map(I => FE_PHN130_framebuffer_buf_92_2380, Z => FE_PHN182_framebuffer_buf_92_2380);
  FE_PHC181_framebuffer_buf_39_2327 : DEL01BWP7T port map(I => FE_PHN173_framebuffer_buf_39_2327, Z => FE_PHN181_framebuffer_buf_39_2327);
  FE_PHC180_framebuffer_buf_105_2393 : DEL01BWP7T port map(I => FE_PHN154_framebuffer_buf_105_2393, Z => FE_PHN180_framebuffer_buf_105_2393);
  FE_PHC179_framebuffer_buf_123_2411 : DEL01BWP7T port map(I => FE_PHN127_framebuffer_buf_123_2411, Z => FE_PHN179_framebuffer_buf_123_2411);
  FE_PHC178_framebuffer_buf_118_2406 : DEL01BWP7T port map(I => FE_PHN149_framebuffer_buf_118_2406, Z => FE_PHN178_framebuffer_buf_118_2406);
  FE_PHC177_framebuffer_buf_151_2439 : DEL01BWP7T port map(I => framebuffer_buf_151_2439, Z => FE_PHN177_framebuffer_buf_151_2439);
  FE_PHC176_calc_buf_out_20_2284 : DEL01BWP7T port map(I => calc_buf_out_20_2284, Z => FE_PHN176_calc_buf_out_20_2284);
  FE_PHC175_framebuffer_buf_109_2397 : DEL3BWP7T port map(I => FE_PHN175_framebuffer_buf_109_2397, Z => framebuffer_buf_109_2397);
  FE_PHC174_framebuffer_buf_20_2308 : BUFFD3BWP7T port map(I => framebuffer_buf_20_2308, Z => FE_PHN174_framebuffer_buf_20_2308);
  FE_PHC173_framebuffer_buf_39_2327 : CKBD2BWP7T port map(I => framebuffer_buf_39_2327, Z => FE_PHN173_framebuffer_buf_39_2327);
  FE_PHC172_framebuffer_buf_134_2422 : BUFFD5BWP7T port map(I => framebuffer_buf_134_2422, Z => FE_PHN172_framebuffer_buf_134_2422);
  FE_PHC171_framebuffer_buf_44_2332 : DEL1BWP7T port map(I => FE_PHN171_framebuffer_buf_44_2332, Z => framebuffer_buf_44_2332);
  FE_PHC170_framebuffer_buf_131_2419 : DEL1BWP7T port map(I => framebuffer_buf_131_2419, Z => FE_PHN170_framebuffer_buf_131_2419);
  FE_PHC169_calc_buf_out_20_2284 : CKBD0BWP7T port map(I => FE_PHN176_calc_buf_out_20_2284, Z => FE_PHN169_calc_buf_out_20_2284);
  FE_PHC168_framebuffer_buf_56_2344 : CKBD3BWP7T port map(I => framebuffer_buf_56_2344, Z => FE_PHN168_framebuffer_buf_56_2344);
  FE_PHC167_framebuffer_buf_130_2418 : DEL1BWP7T port map(I => FE_PHN167_framebuffer_buf_130_2418, Z => framebuffer_buf_130_2418);
  FE_PHC166_framebuffer_buf_1_2289 : DEL0BWP7T port map(I => framebuffer_buf_1_2289, Z => FE_PHN166_framebuffer_buf_1_2289);
  FE_PHC165_framebuffer_buf_50_2338 : CKBD4BWP7T port map(I => framebuffer_buf_50_2338, Z => FE_PHN165_framebuffer_buf_50_2338);
  FE_PHC164_framebuffer_buf_129_2417 : DEL0BWP7T port map(I => framebuffer_buf_129_2417, Z => FE_PHN164_framebuffer_buf_129_2417);
  FE_PHC163_framebuffer_buf_93_2381 : DEL0BWP7T port map(I => framebuffer_buf_93_2381, Z => FE_PHN163_framebuffer_buf_93_2381);
  FE_PHC162_framebuffer_buf_151_2439 : CKBD0BWP7T port map(I => FE_PHN162_framebuffer_buf_151_2439, Z => framebuffer_buf_151_2439);
  FE_PHC161_framebuffer_buf_136_2424 : DEL0BWP7T port map(I => FE_PHN161_framebuffer_buf_136_2424, Z => framebuffer_buf_136_2424);
  FE_PHC160_framebuffer_buf_10_2298 : CKBD0BWP7T port map(I => framebuffer_buf_10_2298, Z => FE_PHN160_framebuffer_buf_10_2298);
  FE_PHC159_framebuffer_buf_150_2438 : CKBD0BWP7T port map(I => FE_PHN159_framebuffer_buf_150_2438, Z => framebuffer_buf_150_2438);
  FE_PHC158_framebuffer_buf_117_2405 : DEL0BWP7T port map(I => framebuffer_buf_117_2405, Z => FE_PHN158_framebuffer_buf_117_2405);
  FE_PHC157_framebuffer_buf_104_2392 : CKBD0BWP7T port map(I => framebuffer_buf_104_2392, Z => FE_PHN157_framebuffer_buf_104_2392);
  FE_PHC156_framebuffer_buf_143_2431 : DEL0BWP7T port map(I => framebuffer_buf_143_2431, Z => FE_PHN156_framebuffer_buf_143_2431);
  FE_PHC155_framebuffer_buf_138_2426 : DEL0BWP7T port map(I => FE_PHN155_framebuffer_buf_138_2426, Z => framebuffer_buf_138_2426);
  FE_PHC154_framebuffer_buf_105_2393 : CKBD0BWP7T port map(I => framebuffer_buf_105_2393, Z => FE_PHN154_framebuffer_buf_105_2393);
  FE_PHC153_framebuffer_buf_108_2396 : DEL0BWP7T port map(I => framebuffer_buf_108_2396, Z => FE_PHN153_framebuffer_buf_108_2396);
  FE_PHC152_framebuffer_buf_43_2331 : CKBD4BWP7T port map(I => framebuffer_buf_43_2331, Z => FE_PHN152_framebuffer_buf_43_2331);
  FE_PHC151_framebuffer_buf_75_2363 : DEL0BWP7T port map(I => framebuffer_buf_75_2363, Z => FE_PHN151_framebuffer_buf_75_2363);
  FE_PHC150_calc_buf_out_21_2285 : DEL0BWP7T port map(I => calc_buf_out_21_2285, Z => FE_PHN150_calc_buf_out_21_2285);
  FE_PHC149_framebuffer_buf_118_2406 : CKBD0BWP7T port map(I => framebuffer_buf_118_2406, Z => FE_PHN149_framebuffer_buf_118_2406);
  FE_PHC148_framebuffer_buf_78_2366 : CKBD3BWP7T port map(I => FE_PHN148_framebuffer_buf_78_2366, Z => framebuffer_buf_78_2366);
  FE_PHC147_framebuffer_buf_32_2320 : CKBD3BWP7T port map(I => FE_PHN147_framebuffer_buf_32_2320, Z => framebuffer_buf_32_2320);
  FE_PHC146_framebuffer_buf_107_2395 : CKBD3BWP7T port map(I => framebuffer_buf_107_2395, Z => FE_PHN146_framebuffer_buf_107_2395);
  FE_PHC145_framebuffer_buf_84_2372 : DEL0BWP7T port map(I => framebuffer_buf_84_2372, Z => FE_PHN145_framebuffer_buf_84_2372);
  FE_PHC144_framebuffer_buf_23_2311 : DEL0BWP7T port map(I => framebuffer_buf_23_2311, Z => FE_PHN144_framebuffer_buf_23_2311);
  FE_PHC143_framebuffer_buf_14_2302 : CKBD0BWP7T port map(I => framebuffer_buf_14_2302, Z => FE_PHN143_framebuffer_buf_14_2302);
  FE_PHC142_framebuffer_buf_62_2350 : DEL0BWP7T port map(I => framebuffer_buf_62_2350, Z => FE_PHN142_framebuffer_buf_62_2350);
  FE_PHC141_calc_buf_out_19_2283 : DEL0BWP7T port map(I => calc_buf_out_19_2283, Z => FE_PHN141_calc_buf_out_19_2283);
  FE_PHC140_framebuffer_buf_42_2330 : DEL0BWP7T port map(I => framebuffer_buf_42_2330, Z => FE_PHN140_framebuffer_buf_42_2330);
  FE_PHC139_framebuffer_buf_153_2441 : CKBD0BWP7T port map(I => framebuffer_buf_153_2441, Z => FE_PHN139_framebuffer_buf_153_2441);
  FE_PHC138_framebuffer_buf_60_2348 : DEL0BWP7T port map(I => framebuffer_buf_60_2348, Z => FE_PHN138_framebuffer_buf_60_2348);
  FE_PHC137_framebuffer_buf_80_2368 : DEL0BWP7T port map(I => framebuffer_buf_80_2368, Z => FE_PHN137_framebuffer_buf_80_2368);
  FE_PHC136_framebuffer_buf_71_2359 : DEL0BWP7T port map(I => framebuffer_buf_71_2359, Z => FE_PHN136_framebuffer_buf_71_2359);
  FE_PHC135_framebuffer_buf_47_2335 : DEL0BWP7T port map(I => FE_PHN135_framebuffer_buf_47_2335, Z => framebuffer_buf_47_2335);
  FE_PHC134_framebuffer_buf_99_2387 : DEL0BWP7T port map(I => FE_PHN134_framebuffer_buf_99_2387, Z => framebuffer_buf_99_2387);
  FE_PHC133_framebuffer_buf_21_2309 : CKBD3BWP7T port map(I => framebuffer_buf_21_2309, Z => FE_PHN133_framebuffer_buf_21_2309);
  FE_PHC132_framebuffer_buf_28_2316 : DEL0BWP7T port map(I => framebuffer_buf_28_2316, Z => FE_PHN132_framebuffer_buf_28_2316);
  FE_PHC131_framebuffer_buf_16_2304 : DEL0BWP7T port map(I => framebuffer_buf_16_2304, Z => FE_PHN131_framebuffer_buf_16_2304);
  FE_PHC130_framebuffer_buf_92_2380 : CKBD0BWP7T port map(I => framebuffer_buf_92_2380, Z => FE_PHN130_framebuffer_buf_92_2380);
  FE_PHC129_framebuffer_buf_26_2314 : DEL0BWP7T port map(I => framebuffer_buf_26_2314, Z => FE_PHN129_framebuffer_buf_26_2314);
  FE_PHC128_framebuffer_buf_29_2317 : DEL0BWP7T port map(I => framebuffer_buf_29_2317, Z => FE_PHN128_framebuffer_buf_29_2317);
  FE_PHC127_framebuffer_buf_123_2411 : CKBD0BWP7T port map(I => framebuffer_buf_123_2411, Z => FE_PHN127_framebuffer_buf_123_2411);
  FE_PHC126_framebuffer_buf_8_2296 : DEL0BWP7T port map(I => framebuffer_buf_8_2296, Z => FE_PHN126_framebuffer_buf_8_2296);
  FE_PHC125_framebuffer_buf_114_2402 : DEL0BWP7T port map(I => framebuffer_buf_114_2402, Z => FE_PHN125_framebuffer_buf_114_2402);
  FE_PHC124_framebuffer_buf_73_2361 : DEL0BWP7T port map(I => framebuffer_buf_73_2361, Z => FE_PHN124_framebuffer_buf_73_2361);
  FE_PHC123_framebuffer_buf_35_2323 : DEL0BWP7T port map(I => framebuffer_buf_35_2323, Z => FE_PHN123_framebuffer_buf_35_2323);
  FE_PHC122_framebuffer_buf_12_2300 : DEL0BWP7T port map(I => FE_PHN122_framebuffer_buf_12_2300, Z => framebuffer_buf_12_2300);
  FE_PHC121_framebuffer_buf_3_2291 : CKBD3BWP7T port map(I => FE_PHN121_framebuffer_buf_3_2291, Z => framebuffer_buf_3_2291);
  FE_PHC120_framebuffer_buf_31_2319 : DEL0BWP7T port map(I => framebuffer_buf_31_2319, Z => FE_PHN120_framebuffer_buf_31_2319);
  FE_PHC119_framebuffer_buf_66_2354 : CKBD0BWP7T port map(I => framebuffer_buf_66_2354, Z => FE_PHN119_framebuffer_buf_66_2354);
  FE_PHC118_framebuffer_buf_154_2442 : CKBD3BWP7T port map(I => framebuffer_buf_154_2442, Z => FE_PHN118_framebuffer_buf_154_2442);
  FE_PHC117_framebuffer_buf_102_2390 : DEL0BWP7T port map(I => framebuffer_buf_102_2390, Z => FE_PHN117_framebuffer_buf_102_2390);
  FE_PHC116_framebuffer_buf_55_2343 : DEL0BWP7T port map(I => framebuffer_buf_55_2343, Z => FE_PHN116_framebuffer_buf_55_2343);
  FE_PHC115_framebuffer_buf_27_2315 : DEL0BWP7T port map(I => framebuffer_buf_27_2315, Z => FE_PHN115_framebuffer_buf_27_2315);
  FE_PHC114_framebuffer_buf_85_2373 : DEL0BWP7T port map(I => framebuffer_buf_85_2373, Z => FE_PHN114_framebuffer_buf_85_2373);
  FE_PHC113_framebuffer_buf_37_2325 : CKBD3BWP7T port map(I => framebuffer_buf_37_2325, Z => FE_PHN113_framebuffer_buf_37_2325);
  FE_PHC112_framebuffer_buf_25_2313 : DEL0BWP7T port map(I => framebuffer_buf_25_2313, Z => FE_PHN112_framebuffer_buf_25_2313);
  FE_PHC111_framebuffer_buf_113_2401 : DEL0BWP7T port map(I => framebuffer_buf_113_2401, Z => FE_PHN111_framebuffer_buf_113_2401);
  FE_PHC110_calc_buf_out_15_2279 : DEL0BWP7T port map(I => calc_buf_out_15_2279, Z => FE_PHN110_calc_buf_out_15_2279);
  FE_PHC109_framebuffer_buf_46_2334 : DEL0BWP7T port map(I => framebuffer_buf_46_2334, Z => FE_PHN109_framebuffer_buf_46_2334);
  FE_PHC108_framebuffer_buf_126_2414 : DEL0BWP7T port map(I => framebuffer_buf_126_2414, Z => FE_PHN108_framebuffer_buf_126_2414);
  FE_PHC107_framebuffer_buf_135_2423 : DEL0BWP7T port map(I => FE_PHN107_framebuffer_buf_135_2423, Z => framebuffer_buf_135_2423);
  FE_PHC106_framebuffer_buf_59_2347 : DEL0BWP7T port map(I => FE_PHN106_framebuffer_buf_59_2347, Z => framebuffer_buf_59_2347);
  FE_PHC105_framebuffer_buf_145_2433 : DEL0BWP7T port map(I => framebuffer_buf_145_2433, Z => FE_PHN105_framebuffer_buf_145_2433);
  FE_PHC104_framebuffer_buf_36_2324 : DEL0BWP7T port map(I => framebuffer_buf_36_2324, Z => FE_PHN104_framebuffer_buf_36_2324);
  FE_PHC103_framebuffer_buf_34_2322 : DEL0BWP7T port map(I => framebuffer_buf_34_2322, Z => FE_PHN103_framebuffer_buf_34_2322);
  FE_PHC102_framebuffer_buf_81_2369 : DEL0BWP7T port map(I => framebuffer_buf_81_2369, Z => FE_PHN102_framebuffer_buf_81_2369);
  FE_PHC101_framebuffer_buf_5_2293 : DEL0BWP7T port map(I => framebuffer_buf_5_2293, Z => FE_PHN101_framebuffer_buf_5_2293);
  FE_PHC100_framebuffer_buf_86_2374 : CKBD3BWP7T port map(I => framebuffer_buf_86_2374, Z => FE_PHN100_framebuffer_buf_86_2374);
  FE_PHC99_framebuffer_buf_137_2425 : DEL0BWP7T port map(I => FE_PHN99_framebuffer_buf_137_2425, Z => framebuffer_buf_137_2425);
  FE_PHC98_framebuffer_buf_98_2386 : DEL0BWP7T port map(I => FE_PHN98_framebuffer_buf_98_2386, Z => framebuffer_buf_98_2386);
  FE_PHC97_framebuffer_buf_156_2444 : DEL0BWP7T port map(I => framebuffer_buf_156_2444, Z => FE_PHN97_framebuffer_buf_156_2444);
  FE_PHC96_framebuffer_buf_124_2412 : DEL0BWP7T port map(I => framebuffer_buf_124_2412, Z => FE_PHN96_framebuffer_buf_124_2412);
  FE_PHC95_framebuffer_buf_38_2326 : DEL0BWP7T port map(I => framebuffer_buf_38_2326, Z => FE_PHN95_framebuffer_buf_38_2326);
  FE_PHC94_framebuffer_buf_140_2428 : DEL0BWP7T port map(I => framebuffer_buf_140_2428, Z => FE_PHN94_framebuffer_buf_140_2428);
  FE_PHC93_calc_buf_out_12_2276 : DEL0BWP7T port map(I => FE_PHN93_calc_buf_out_12_2276, Z => calc_buf_out_12_2276);
  FE_PHC92_framebuffer_buf_7_2295 : CKBD3BWP7T port map(I => framebuffer_buf_7_2295, Z => FE_PHN92_framebuffer_buf_7_2295);
  FE_PHC91_framebuffer_buf_132_2420 : DEL0BWP7T port map(I => framebuffer_buf_132_2420, Z => FE_PHN91_framebuffer_buf_132_2420);
  FE_PHC90_framebuffer_buf_45_2333 : DEL0BWP7T port map(I => framebuffer_buf_45_2333, Z => FE_PHN90_framebuffer_buf_45_2333);
  FE_PHC89_framebuffer_buf_88_2376 : CKBD3BWP7T port map(I => framebuffer_buf_88_2376, Z => FE_PHN89_framebuffer_buf_88_2376);
  FE_PHC88_framebuffer_buf_139_2427 : DEL0BWP7T port map(I => FE_PHN88_framebuffer_buf_139_2427, Z => framebuffer_buf_139_2427);
  FE_PHC87_framebuffer_buf_142_2430 : DEL0BWP7T port map(I => FE_PHN87_framebuffer_buf_142_2430, Z => framebuffer_buf_142_2430);
  FE_PHC86_framebuffer_buf_54_2342 : CKBD3BWP7T port map(I => framebuffer_buf_54_2342, Z => FE_PHN86_framebuffer_buf_54_2342);
  FE_PHC85_framebuffer_buf_48_2336 : DEL0BWP7T port map(I => framebuffer_buf_48_2336, Z => FE_PHN85_framebuffer_buf_48_2336);
  FE_PHC84_framebuffer_buf_70_2358 : DEL0BWP7T port map(I => framebuffer_buf_70_2358, Z => FE_PHN84_framebuffer_buf_70_2358);
  FE_PHC83_framebuffer_buf_33_2321 : DEL0BWP7T port map(I => framebuffer_buf_33_2321, Z => FE_PHN83_framebuffer_buf_33_2321);
  FE_PHC82_framebuffer_buf_24_2312 : DEL0BWP7T port map(I => framebuffer_buf_24_2312, Z => FE_PHN82_framebuffer_buf_24_2312);
  FE_PHC81_framebuffer_buf_76_2364 : CKBD3BWP7T port map(I => framebuffer_buf_76_2364, Z => FE_PHN81_framebuffer_buf_76_2364);
  FE_PHC80_framebuffer_buf_146_2434 : DEL0BWP7T port map(I => framebuffer_buf_146_2434, Z => FE_PHN80_framebuffer_buf_146_2434);
  FE_PHC79_framebuffer_buf_91_2379 : DEL0BWP7T port map(I => framebuffer_buf_91_2379, Z => FE_PHN79_framebuffer_buf_91_2379);
  FE_PHC78_framebuffer_buf_63_2351 : DEL0BWP7T port map(I => framebuffer_buf_63_2351, Z => FE_PHN78_framebuffer_buf_63_2351);
  FE_PHC77_framebuffer_buf_17_2305 : DEL0BWP7T port map(I => framebuffer_buf_17_2305, Z => FE_PHN77_framebuffer_buf_17_2305);
  FE_PHC76_framebuffer_buf_30_2318 : DEL0BWP7T port map(I => framebuffer_buf_30_2318, Z => FE_PHN76_framebuffer_buf_30_2318);
  FE_PHC75_framebuffer_buf_120_2408 : DEL0BWP7T port map(I => framebuffer_buf_120_2408, Z => FE_PHN75_framebuffer_buf_120_2408);
  FE_PHC74_framebuffer_buf_116_2404 : DEL0BWP7T port map(I => framebuffer_buf_116_2404, Z => FE_PHN74_framebuffer_buf_116_2404);
  FE_PHC73_framebuffer_buf_52_2340 : DEL0BWP7T port map(I => framebuffer_buf_52_2340, Z => FE_PHN73_framebuffer_buf_52_2340);
  FE_PHC72_framebuffer_buf_87_2375 : DEL0BWP7T port map(I => framebuffer_buf_87_2375, Z => FE_PHN72_framebuffer_buf_87_2375);
  FE_PHC71_framebuffer_buf_111_2399 : DEL0BWP7T port map(I => framebuffer_buf_111_2399, Z => FE_PHN71_framebuffer_buf_111_2399);
  FE_PHC70_framebuffer_buf_100_2388 : DEL0BWP7T port map(I => framebuffer_buf_100_2388, Z => FE_PHN70_framebuffer_buf_100_2388);
  FE_PHC69_framebuffer_buf_2_2290 : DEL0BWP7T port map(I => framebuffer_buf_2_2290, Z => FE_PHN69_framebuffer_buf_2_2290);
  FE_PHC68_framebuffer_buf_9_2297 : DEL0BWP7T port map(I => framebuffer_buf_9_2297, Z => FE_PHN68_framebuffer_buf_9_2297);
  FE_PHC67_framebuffer_buf_6_2294 : DEL0BWP7T port map(I => framebuffer_buf_6_2294, Z => FE_PHN67_framebuffer_buf_6_2294);
  FE_PHC66_framebuffer_buf_41_2329 : DEL0BWP7T port map(I => framebuffer_buf_41_2329, Z => FE_PHN66_framebuffer_buf_41_2329);
  FE_PHC65_framebuffer_buf_125_2413 : DEL0BWP7T port map(I => framebuffer_buf_125_2413, Z => FE_PHN65_framebuffer_buf_125_2413);
  FE_PHC64_framebuffer_buf_64_2352 : DEL0BWP7T port map(I => framebuffer_buf_64_2352, Z => FE_PHN64_framebuffer_buf_64_2352);
  FE_PHC63_framebuffer_buf_95_2383 : DEL0BWP7T port map(I => framebuffer_buf_95_2383, Z => FE_PHN63_framebuffer_buf_95_2383);
  FE_PHC62_framebuffer_buf_94_2382 : DEL0BWP7T port map(I => framebuffer_buf_94_2382, Z => FE_PHN62_framebuffer_buf_94_2382);
  FE_PHC61_calc_buf_out_23_2287 : DEL0BWP7T port map(I => calc_buf_out_23_2287, Z => FE_PHN61_calc_buf_out_23_2287);
  FE_PHC60_framebuffer_buf_0_2288 : DEL0BWP7T port map(I => framebuffer_buf_0_2288, Z => FE_PHN60_framebuffer_buf_0_2288);
  FE_PHC59_framebuffer_buf_112_2400 : DEL0BWP7T port map(I => framebuffer_buf_112_2400, Z => FE_PHN59_framebuffer_buf_112_2400);
  FE_PHC58_framebuffer_buf_51_2339 : DEL0BWP7T port map(I => framebuffer_buf_51_2339, Z => FE_PHN58_framebuffer_buf_51_2339);
  FE_PHC57_framebuffer_buf_58_2346 : DEL0BWP7T port map(I => framebuffer_buf_58_2346, Z => FE_PHN57_framebuffer_buf_58_2346);
  FE_PHC56_framebuffer_buf_103_2391 : DEL0BWP7T port map(I => framebuffer_buf_103_2391, Z => FE_PHN56_framebuffer_buf_103_2391);
  FE_PHC55_framebuffer_buf_101_2389 : DEL0BWP7T port map(I => framebuffer_buf_101_2389, Z => FE_PHN55_framebuffer_buf_101_2389);
  FE_PHC54_framebuffer_buf_96_2384 : DEL0BWP7T port map(I => framebuffer_buf_96_2384, Z => FE_PHN54_framebuffer_buf_96_2384);
  FE_PHC53_framebuffer_buf_69_2357 : BUFFD3BWP7T port map(I => framebuffer_buf_69_2357, Z => FE_PHN53_framebuffer_buf_69_2357);
  FE_PHC52_framebuffer_buf_110_2398 : DEL0BWP7T port map(I => framebuffer_buf_110_2398, Z => FE_PHN52_framebuffer_buf_110_2398);
  FE_PHC51_framebuffer_buf_128_2416 : DEL0BWP7T port map(I => FE_PHN51_framebuffer_buf_128_2416, Z => framebuffer_buf_128_2416);
  FE_PHC50_framebuffer_buf_4_2292 : DEL0BWP7T port map(I => FE_PHN50_framebuffer_buf_4_2292, Z => framebuffer_buf_4_2292);
  FE_PHC49_framebuffer_buf_141_2429 : CKBD3BWP7T port map(I => framebuffer_buf_141_2429, Z => FE_PHN49_framebuffer_buf_141_2429);
  FE_PHC48_framebuffer_buf_72_2360 : DEL0BWP7T port map(I => framebuffer_buf_72_2360, Z => FE_PHN48_framebuffer_buf_72_2360);
  FE_PHC47_framebuffer_buf_106_2394 : DEL0BWP7T port map(I => framebuffer_buf_106_2394, Z => FE_PHN47_framebuffer_buf_106_2394);
  FE_PHC46_framebuffer_buf_97_2385 : DEL0BWP7T port map(I => framebuffer_buf_97_2385, Z => FE_PHN46_framebuffer_buf_97_2385);
  FE_PHC45_framebuffer_buf_122_2410 : BUFFD3BWP7T port map(I => framebuffer_buf_122_2410, Z => FE_PHN45_framebuffer_buf_122_2410);
  FE_PHC44_framebuffer_buf_157_2445 : BUFFD3BWP7T port map(I => framebuffer_buf_157_2445, Z => FE_PHN44_framebuffer_buf_157_2445);
  FE_PHC43_framebuffer_buf_53_2341 : BUFFD3BWP7T port map(I => framebuffer_buf_53_2341, Z => FE_PHN43_framebuffer_buf_53_2341);
  FE_PHC42_framebuffer_buf_19_2307 : BUFFD3BWP7T port map(I => framebuffer_buf_19_2307, Z => FE_PHN42_framebuffer_buf_19_2307);
  FE_PHC41_calc_buf_out_16_2280 : DEL0BWP7T port map(I => FE_PHN41_calc_buf_out_16_2280, Z => calc_buf_out_16_2280);
  FE_PHC40_framebuffer_buf_61_2349 : BUFFD3BWP7T port map(I => framebuffer_buf_61_2349, Z => FE_PHN40_framebuffer_buf_61_2349);
  FE_PHC39_calc_buf_out_10_2274 : DEL0BWP7T port map(I => calc_buf_out_10_2274, Z => FE_PHN39_calc_buf_out_10_2274);
  FE_PHC38_framebuffer_buf_144_2432 : BUFFD3BWP7T port map(I => framebuffer_buf_144_2432, Z => FE_PHN38_framebuffer_buf_144_2432);
  FE_PHC37_calc_buf_out_13_2277 : DEL0BWP7T port map(I => FE_PHN37_calc_buf_out_13_2277, Z => calc_buf_out_13_2277);
  FE_PHC36_framebuffer_buf_119_2407 : BUFFD3BWP7T port map(I => framebuffer_buf_119_2407, Z => FE_PHN36_framebuffer_buf_119_2407);
  FE_PHC35_calc_buf_out_9_2273 : DEL0BWP7T port map(I => calc_buf_out_9_2273, Z => FE_PHN35_calc_buf_out_9_2273);
  FE_PHC34_framebuffer_buf_68_2356 : BUFFD3BWP7T port map(I => framebuffer_buf_68_2356, Z => FE_PHN34_framebuffer_buf_68_2356);
  FE_PHC33_framebuffer_buf_11_2299 : BUFFD3BWP7T port map(I => framebuffer_buf_11_2299, Z => FE_PHN33_framebuffer_buf_11_2299);
  FE_PHC32_calc_buf_out_14_2278 : DEL0BWP7T port map(I => calc_buf_out_14_2278, Z => FE_PHN32_calc_buf_out_14_2278);
  FE_PHC31_framebuffer_buf_89_2377 : BUFFD3BWP7T port map(I => framebuffer_buf_89_2377, Z => FE_PHN31_framebuffer_buf_89_2377);
  FE_PHC30_framebuffer_buf_18_2306 : BUFFD3BWP7T port map(I => framebuffer_buf_18_2306, Z => FE_PHN30_framebuffer_buf_18_2306);
  FE_PHC29_framebuffer_buf_121_2409 : BUFFD3BWP7T port map(I => framebuffer_buf_121_2409, Z => FE_PHN29_framebuffer_buf_121_2409);
  FE_PHC28_calc_buf_out_22_2286 : DEL0BWP7T port map(I => FE_PHN28_calc_buf_out_22_2286, Z => calc_buf_out_22_2286);
  FE_PHC27_framebuffer_buf_127_2415 : BUFFD3BWP7T port map(I => framebuffer_buf_127_2415, Z => FE_PHN27_framebuffer_buf_127_2415);
  FE_PHC26_calc_buf_out_18_2282 : DEL0BWP7T port map(I => calc_buf_out_18_2282, Z => FE_PHN26_calc_buf_out_18_2282);
  FE_PHC25_calc_buf_out_11_2275 : DEL0BWP7T port map(I => calc_buf_out_11_2275, Z => FE_PHN25_calc_buf_out_11_2275);
  FE_PHC24_framebuffer_buf_155_2443 : BUFFD3BWP7T port map(I => framebuffer_buf_155_2443, Z => FE_PHN24_framebuffer_buf_155_2443);
  FE_PHC23_calc_buf_out_17_2281 : DEL0BWP7T port map(I => FE_PHN23_calc_buf_out_17_2281, Z => calc_buf_out_17_2281);
  FE_PHC22_calc_buf_out_8_2272 : DEL0BWP7T port map(I => calc_buf_out_8_2272, Z => FE_PHN22_calc_buf_out_8_2272);
  FE_PHC21_framebuffer_buf_149_2437 : DEL01BWP7T port map(I => framebuffer_buf_149_2437, Z => FE_PHN21_framebuffer_buf_149_2437);
  FE_PHC20_framebuffer_buf_79_2367 : CKBD0BWP7T port map(I => framebuffer_buf_79_2367, Z => FE_PHN20_framebuffer_buf_79_2367);
  FE_PHC19_framebuffer_buf_15_2303 : DEL01BWP7T port map(I => framebuffer_buf_15_2303, Z => FE_PHN19_framebuffer_buf_15_2303);
  FE_PHC18_framebuffer_buf_22_2310 : CKBD0BWP7T port map(I => framebuffer_buf_22_2310, Z => FE_PHN18_framebuffer_buf_22_2310);
  FE_PHC17_framebuffer_buf_74_2362 : CKBD0BWP7T port map(I => framebuffer_buf_74_2362, Z => FE_PHN17_framebuffer_buf_74_2362);
  FE_PHC16_framebuffer_buf_65_2353 : CKBD0BWP7T port map(I => framebuffer_buf_65_2353, Z => FE_PHN16_framebuffer_buf_65_2353);
  FE_PHC15_framebuffer_buf_77_2365 : CKBD0BWP7T port map(I => framebuffer_buf_77_2365, Z => FE_PHN15_framebuffer_buf_77_2365);
  FE_PHC14_framebuffer_buf_13_2301 : CKBD0BWP7T port map(I => framebuffer_buf_13_2301, Z => FE_PHN14_framebuffer_buf_13_2301);
  FE_PHC13_framebuffer_buf_148_2436 : CKBD0BWP7T port map(I => framebuffer_buf_148_2436, Z => FE_PHN13_framebuffer_buf_148_2436);
  FE_PHC12_framebuffer_buf_67_2355 : CKBD0BWP7T port map(I => framebuffer_buf_67_2355, Z => FE_PHN12_framebuffer_buf_67_2355);
  FE_PHC11_framebuffer_buf_57_2345 : CKBD0BWP7T port map(I => framebuffer_buf_57_2345, Z => FE_PHN11_framebuffer_buf_57_2345);
  FE_PHC10_framebuffer_buf_83_2371 : CKBD0BWP7T port map(I => framebuffer_buf_83_2371, Z => FE_PHN10_framebuffer_buf_83_2371);
  FE_PHC9_framebuffer_buf_90_2378 : CKBD0BWP7T port map(I => framebuffer_buf_90_2378, Z => FE_PHN9_framebuffer_buf_90_2378);
  FE_PHC8_framebuffer_buf_49_2337 : CKBD0BWP7T port map(I => framebuffer_buf_49_2337, Z => FE_PHN8_framebuffer_buf_49_2337);
  FE_PHC7_framebuffer_buf_152_2440 : CKBD0BWP7T port map(I => framebuffer_buf_152_2440, Z => FE_PHN7_framebuffer_buf_152_2440);
  FE_PHC6_framebuffer_buf_133_2421 : CKBD0BWP7T port map(I => framebuffer_buf_133_2421, Z => FE_PHN6_framebuffer_buf_133_2421);
  FE_PHC5_framebuffer_buf_82_2370 : CKBD0BWP7T port map(I => FE_PHN5_framebuffer_buf_82_2370, Z => framebuffer_buf_82_2370);
  FE_PHC4_framebuffer_buf_115_2403 : CKBD0BWP7T port map(I => framebuffer_buf_115_2403, Z => FE_PHN4_framebuffer_buf_115_2403);
  FE_PHC3_framebuffer_buf_40_2328 : CKBD0BWP7T port map(I => framebuffer_buf_40_2328, Z => FE_PHN3_framebuffer_buf_40_2328);
  FE_PHC2_framebuffer_buf_147_2435 : CKBD0BWP7T port map(I => framebuffer_buf_147_2435, Z => FE_PHN2_framebuffer_buf_147_2435);
  FE_OFC1_FE_DBTN0_reset : BUFFD2BWP7T port map(I => FE_OFN0_FE_DBTN0_reset, Z => FE_OFN1_FE_DBTN0_reset);
  FE_OFC0_FE_DBTN0_reset : BUFFD2BWP7T port map(I => FE_DBTN0_reset, Z => FE_OFN0_FE_DBTN0_reset);
  CTS_ccl_a_BUF_clk_G0_L2_2 : CKBD12BWP7T port map(I => CTS_14, Z => CTS_13);
  CTS_ccl_a_BUF_clk_G0_L2_1 : CKBD12BWP7T port map(I => CTS_14, Z => CTS_12);
  CTS_ccl_a_BUF_clk_G0_L1_1 : CKBD6BWP7T port map(I => clk, Z => CTS_14);
  FE_DBTC0_reset : INVD2BWP7T port map(I => reset, ZN => FE_DBTN0_reset);
  counter_reg_6 : DFKCNQD1BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => new_counter(6), Q => counter(6));
  new_counter_reg_7 : LHQD1BWP7T port map(D => n_395, E => n_396, Q => new_counter(7));
  new_calc_buf_out_reg_1 : LHQD1BWP7T port map(D => n_372, E => n_397, Q => new_calc_buf_out(1));
  new_calc_buf_out_reg_5 : LHQD1BWP7T port map(D => n_393, E => n_397, Q => new_calc_buf_out(5));
  new_calc_buf_out_reg_3 : LHQD1BWP7T port map(D => n_388, E => n_397, Q => new_calc_buf_out(3));
  new_calc_buf_out_reg_2 : LHQD1BWP7T port map(D => n_356, E => n_397, Q => new_calc_buf_out(2));
  new_calc_buf_out_reg_4 : LHQD1BWP7T port map(D => n_373, E => n_397, Q => new_calc_buf_out(4));
  new_calc_buf_out_reg_0 : LHQD1BWP7T port map(D => n_357, E => n_397, Q => new_calc_buf_out(0));
  new_calc_buf_out_reg_7 : LHQD1BWP7T port map(D => n_389, E => n_397, Q => new_calc_buf_out(7));
  new_calc_buf_out_reg_6 : LHQD1BWP7T port map(D => n_392, E => n_397, Q => new_calc_buf_out(6));
  new_counter_reg_0 : LHQD1BWP7T port map(D => n_327, E => n_396, Q => new_counter(0));
  new_counter_reg_6 : LHQD1BWP7T port map(D => n_311, E => n_396, Q => new_counter(6));
  g23098 : AO32D0BWP7T port map(A1 => n_99, A2 => counter(5), A3 => counter(6), B1 => n_156, B2 => counter(7), Z => n_395);
  g23330 : AO22D0BWP7T port map(A1 => n_377, A2 => FE_PHN141_calc_buf_out_19_2283, B1 => sqi_data_in(3), B2 => n_376, Z => n_394);
  g23312 : AO22D0BWP7T port map(A1 => n_391, A2 => calc_buf_out_5_2269, B1 => sqi_data_in(5), B2 => n_390, Z => n_393);
  g23313 : AO22D0BWP7T port map(A1 => n_391, A2 => calc_buf_out_6_2270, B1 => sqi_data_in(6), B2 => n_390, Z => n_392);
  g23314 : AO22D0BWP7T port map(A1 => n_391, A2 => calc_buf_out_7_2271, B1 => sqi_data_in(7), B2 => n_390, Z => n_389);
  g23316 : AO22D0BWP7T port map(A1 => n_391, A2 => calc_buf_out_3_2267, B1 => sqi_data_in(3), B2 => n_390, Z => n_388);
  g23320 : AO22D0BWP7T port map(A1 => n_385, A2 => FE_PHN22_calc_buf_out_8_2272, B1 => sqi_data_in(0), B2 => n_384, Z => n_387);
  g23321 : AO22D0BWP7T port map(A1 => n_385, A2 => FE_PHN35_calc_buf_out_9_2273, B1 => sqi_data_in(1), B2 => n_384, Z => n_386);
  g23322 : AO22D0BWP7T port map(A1 => n_385, A2 => FE_PHN39_calc_buf_out_10_2274, B1 => sqi_data_in(2), B2 => n_384, Z => n_383);
  g23323 : AO22D0BWP7T port map(A1 => n_385, A2 => FE_PHN25_calc_buf_out_11_2275, B1 => sqi_data_in(3), B2 => n_384, Z => n_382);
  g23324 : AO22D0BWP7T port map(A1 => n_385, A2 => calc_buf_out_12_2276, B1 => sqi_data_in(4), B2 => n_384, Z => n_381);
  g23325 : AO22D0BWP7T port map(A1 => n_385, A2 => FE_PHN32_calc_buf_out_14_2278, B1 => sqi_data_in(6), B2 => n_384, Z => n_380);
  g23326 : AO22D0BWP7T port map(A1 => n_385, A2 => FE_PHN110_calc_buf_out_15_2279, B1 => sqi_data_in(7), B2 => n_384, Z => n_379);
  g23327 : AO22D0BWP7T port map(A1 => n_377, A2 => calc_buf_out_16_2280, B1 => sqi_data_in(0), B2 => n_376, Z => n_378);
  g23328 : AO22D0BWP7T port map(A1 => n_377, A2 => calc_buf_out_17_2281, B1 => sqi_data_in(1), B2 => n_376, Z => n_375);
  g23329 : AO22D0BWP7T port map(A1 => n_377, A2 => FE_PHN26_calc_buf_out_18_2282, B1 => sqi_data_in(2), B2 => n_376, Z => n_374);
  g23311 : AO22D0BWP7T port map(A1 => n_391, A2 => calc_buf_out_4_2268, B1 => sqi_data_in(4), B2 => n_390, Z => n_373);
  g23306 : AO22D0BWP7T port map(A1 => n_391, A2 => calc_buf_out_1_2265, B1 => sqi_data_in(1), B2 => n_390, Z => n_372);
  g23429 : MOAI22D0BWP7T port map(A1 => n_1522, A2 => n_353, B1 => n_366, B2 => framebuffer_buf_136_2424, ZN => n_371);
  g23332 : AO22D0BWP7T port map(A1 => n_377, A2 => FE_PHN150_calc_buf_out_21_2285, B1 => sqi_data_in(5), B2 => n_376, Z => n_370);
  g23333 : AO22D0BWP7T port map(A1 => n_377, A2 => calc_buf_out_22_2286, B1 => sqi_data_in(6), B2 => n_376, Z => n_369);
  g23432 : MOAI22D0BWP7T port map(A1 => n_1522, A2 => n_350, B1 => n_366, B2 => framebuffer_buf_137_2425, ZN => n_368);
  g23334 : AO22D0BWP7T port map(A1 => n_377, A2 => FE_PHN61_calc_buf_out_23_2287, B1 => sqi_data_in(7), B2 => n_376, Z => n_365);
  g23433 : MOAI22D0BWP7T port map(A1 => n_1522, A2 => n_347, B1 => n_366, B2 => framebuffer_buf_138_2426, ZN => n_364);
  g23435 : MOAI22D0BWP7T port map(A1 => n_1522, A2 => n_345, B1 => n_366, B2 => framebuffer_buf_139_2427, ZN => n_363);
  g23335 : AO22D0BWP7T port map(A1 => n_385, A2 => calc_buf_out_13_2277, B1 => sqi_data_in(5), B2 => n_384, Z => n_362);
  g23436 : MOAI22D0BWP7T port map(A1 => n_1522, A2 => n_343, B1 => n_366, B2 => FE_PHN94_framebuffer_buf_140_2428, ZN => n_361);
  g23437 : MOAI22D0BWP7T port map(A1 => n_1522, A2 => n_341, B1 => n_366, B2 => FE_PHN49_framebuffer_buf_141_2429, ZN => n_360);
  g23438 : MOAI22D0BWP7T port map(A1 => n_1522, A2 => n_339, B1 => n_366, B2 => framebuffer_buf_142_2430, ZN => n_359);
  g23439 : MOAI22D0BWP7T port map(A1 => n_1522, A2 => n_336, B1 => n_366, B2 => FE_PHN156_framebuffer_buf_143_2431, ZN => n_358);
  g23304 : AO22D0BWP7T port map(A1 => n_391, A2 => calc_buf_out_0_2264, B1 => sqi_data_in(0), B2 => n_390, Z => n_357);
  g23305 : AO22D0BWP7T port map(A1 => n_391, A2 => calc_buf_out_2_2266, B1 => sqi_data_in(2), B2 => n_390, Z => n_356);
  g23331 : AO22D0BWP7T port map(A1 => n_377, A2 => FE_PHN169_calc_buf_out_20_2284, B1 => sqi_data_in(4), B2 => n_376, Z => n_355);
  g23382 : MOAI22D0BWP7T port map(A1 => n_351, A2 => n_353, B1 => n_349, B2 => FE_PHN126_framebuffer_buf_8_2296, ZN => n_354);
  g23383 : MOAI22D0BWP7T port map(A1 => n_351, A2 => n_350, B1 => n_349, B2 => FE_PHN68_framebuffer_buf_9_2297, ZN => n_352);
  g23384 : MOAI22D0BWP7T port map(A1 => n_351, A2 => n_347, B1 => n_349, B2 => FE_PHN188_framebuffer_buf_10_2298, ZN => n_348);
  g23385 : MOAI22D0BWP7T port map(A1 => n_351, A2 => n_345, B1 => n_349, B2 => FE_PHN33_framebuffer_buf_11_2299, ZN => n_346);
  g23386 : MOAI22D0BWP7T port map(A1 => n_351, A2 => n_343, B1 => n_349, B2 => framebuffer_buf_12_2300, ZN => n_344);
  g23387 : MOAI22D0BWP7T port map(A1 => n_351, A2 => n_341, B1 => n_349, B2 => FE_PHN14_framebuffer_buf_13_2301, ZN => n_342);
  g23388 : MOAI22D0BWP7T port map(A1 => n_337, A2 => n_339, B1 => n_335, B2 => FE_PHN108_framebuffer_buf_126_2414, ZN => n_340);
  g23389 : MOAI22D0BWP7T port map(A1 => n_337, A2 => n_336, B1 => n_335, B2 => FE_PHN27_framebuffer_buf_127_2415, ZN => n_338);
  g23390 : MOAI22D0BWP7T port map(A1 => n_351, A2 => n_339, B1 => n_349, B2 => FE_PHN143_framebuffer_buf_14_2302, ZN => n_334);
  g23391 : MOAI22D0BWP7T port map(A1 => n_351, A2 => n_336, B1 => n_349, B2 => FE_PHN19_framebuffer_buf_15_2303, ZN => n_333);
  g23392 : MOAI22D0BWP7T port map(A1 => n_330, A2 => n_341, B1 => n_329, B2 => FE_PHN113_framebuffer_buf_37_2325, ZN => n_332);
  g23393 : MOAI22D0BWP7T port map(A1 => n_330, A2 => n_353, B1 => n_329, B2 => framebuffer_buf_32_2320, ZN => n_331);
  g23394 : MOAI22D0BWP7T port map(A1 => n_330, A2 => n_350, B1 => n_329, B2 => FE_PHN83_framebuffer_buf_33_2321, ZN => n_328);
  g23315 : MOAI22D0BWP7T port map(A1 => n_122, A2 => counter(0), B1 => n_151, B2 => counter(0), ZN => n_327);
  g23395 : MOAI22D0BWP7T port map(A1 => n_330, A2 => n_347, B1 => n_329, B2 => FE_PHN103_framebuffer_buf_34_2322, ZN => n_326);
  g23396 : MOAI22D0BWP7T port map(A1 => n_330, A2 => n_343, B1 => n_329, B2 => FE_PHN104_framebuffer_buf_36_2324, ZN => n_325);
  g23397 : MOAI22D0BWP7T port map(A1 => n_330, A2 => n_345, B1 => n_329, B2 => FE_PHN123_framebuffer_buf_35_2323, ZN => n_324);
  g23317 : MOAI22D0BWP7T port map(A1 => n_276, A2 => n_336, B1 => n_275, B2 => framebuffer_buf_135_2423, ZN => n_323);
  g23398 : MOAI22D0BWP7T port map(A1 => n_330, A2 => n_339, B1 => n_329, B2 => FE_PHN95_framebuffer_buf_38_2326, ZN => n_322);
  g23399 : MOAI22D0BWP7T port map(A1 => n_330, A2 => n_336, B1 => n_329, B2 => FE_PHN181_framebuffer_buf_39_2327, ZN => n_321);
  g23400 : MOAI22D0BWP7T port map(A1 => n_318, A2 => n_353, B1 => n_317, B2 => FE_PHN85_framebuffer_buf_48_2336, ZN => n_320);
  g23401 : MOAI22D0BWP7T port map(A1 => n_318, A2 => n_350, B1 => n_317, B2 => FE_PHN8_framebuffer_buf_49_2337, ZN => n_319);
  g23318 : MOAI22D0BWP7T port map(A1 => n_318, A2 => n_343, B1 => n_317, B2 => FE_PHN73_framebuffer_buf_52_2340, ZN => n_316);
  g23319 : MOAI22D0BWP7T port map(A1 => n_318, A2 => n_345, B1 => n_317, B2 => FE_PHN58_framebuffer_buf_51_2339, ZN => n_315);
  g23405 : MOAI22D0BWP7T port map(A1 => n_262, A2 => n_343, B1 => n_261, B2 => FE_PHN34_framebuffer_buf_68_2356, ZN => n_314);
  g23406 : MOAI22D0BWP7T port map(A1 => n_318, A2 => n_339, B1 => n_317, B2 => FE_PHN86_framebuffer_buf_54_2342, ZN => n_313);
  g23348 : MOAI22D0BWP7T port map(A1 => n_233, A2 => n_353, B1 => n_232, B2 => FE_PHN3_framebuffer_buf_40_2328, ZN => n_312);
  g23100 : OAI31D0BWP7T port map(A1 => counter(6), A2 => n_145, A3 => n_144, B => n_155, ZN => n_311);
  g23407 : MOAI22D0BWP7T port map(A1 => n_318, A2 => n_336, B1 => n_317, B2 => FE_PHN116_framebuffer_buf_55_2343, ZN => n_310);
  g23408 : MOAI22D0BWP7T port map(A1 => n_1523, A2 => n_353, B1 => n_303, B2 => FE_PHN59_framebuffer_buf_112_2400, ZN => n_309);
  g23462 : MOAI22D0BWP7T port map(A1 => n_225, A2 => n_353, B1 => n_224, B2 => FE_PHN137_framebuffer_buf_80_2368, ZN => n_308);
  g23460 : MOAI22D0BWP7T port map(A1 => n_246, A2 => n_339, B1 => n_245, B2 => framebuffer_buf_78_2366, ZN => n_307);
  g23409 : MOAI22D0BWP7T port map(A1 => n_301, A2 => n_350, B1 => n_300, B2 => FE_PHN77_framebuffer_buf_17_2305, ZN => n_306);
  g23410 : MOAI22D0BWP7T port map(A1 => n_1523, A2 => n_350, B1 => n_303, B2 => FE_PHN111_framebuffer_buf_113_2401, ZN => n_305);
  g23411 : MOAI22D0BWP7T port map(A1 => n_301, A2 => n_347, B1 => n_300, B2 => FE_PHN30_framebuffer_buf_18_2306, ZN => n_302);
  g23412 : MOAI22D0BWP7T port map(A1 => n_1523, A2 => n_347, B1 => n_303, B2 => FE_PHN125_framebuffer_buf_114_2402, ZN => n_299);
  g23413 : MOAI22D0BWP7T port map(A1 => n_1523, A2 => n_345, B1 => n_303, B2 => FE_PHN4_framebuffer_buf_115_2403, ZN => n_298);
  g23414 : MOAI22D0BWP7T port map(A1 => n_1523, A2 => n_343, B1 => n_303, B2 => FE_PHN74_framebuffer_buf_116_2404, ZN => n_297);
  g23415 : MOAI22D0BWP7T port map(A1 => n_301, A2 => n_345, B1 => n_300, B2 => FE_PHN42_framebuffer_buf_19_2307, ZN => n_296);
  g23416 : MOAI22D0BWP7T port map(A1 => n_271, A2 => n_345, B1 => n_270, B2 => FE_PHN24_framebuffer_buf_155_2443, ZN => n_295);
  g23417 : MOAI22D0BWP7T port map(A1 => n_301, A2 => n_343, B1 => n_300, B2 => FE_PHN174_framebuffer_buf_20_2308, ZN => n_294);
  g23418 : MOAI22D0BWP7T port map(A1 => n_1523, A2 => n_341, B1 => n_303, B2 => FE_PHN158_framebuffer_buf_117_2405, ZN => n_293);
  g23419 : MOAI22D0BWP7T port map(A1 => n_1523, A2 => n_339, B1 => n_303, B2 => FE_PHN178_framebuffer_buf_118_2406, ZN => n_292);
  g23420 : MOAI22D0BWP7T port map(A1 => n_1523, A2 => n_336, B1 => n_303, B2 => FE_PHN36_framebuffer_buf_119_2407, ZN => n_291);
  g23421 : MOAI22D0BWP7T port map(A1 => n_301, A2 => n_341, B1 => n_300, B2 => FE_PHN133_framebuffer_buf_21_2309, ZN => n_290);
  g23422 : MOAI22D0BWP7T port map(A1 => n_301, A2 => n_339, B1 => n_300, B2 => FE_PHN18_framebuffer_buf_22_2310, ZN => n_289);
  g23423 : MOAI22D0BWP7T port map(A1 => n_301, A2 => n_336, B1 => n_300, B2 => FE_PHN144_framebuffer_buf_23_2311, ZN => n_288);
  g23424 : MOAI22D0BWP7T port map(A1 => n_285, A2 => n_353, B1 => n_284, B2 => FE_PHN82_framebuffer_buf_24_2312, ZN => n_287);
  g23425 : MOAI22D0BWP7T port map(A1 => n_285, A2 => n_350, B1 => n_284, B2 => FE_PHN112_framebuffer_buf_25_2313, ZN => n_286);
  g23426 : MOAI22D0BWP7T port map(A1 => n_285, A2 => n_347, B1 => n_284, B2 => FE_PHN129_framebuffer_buf_26_2314, ZN => n_283);
  g23427 : MOAI22D0BWP7T port map(A1 => n_285, A2 => n_345, B1 => n_284, B2 => FE_PHN115_framebuffer_buf_27_2315, ZN => n_282);
  g23428 : MOAI22D0BWP7T port map(A1 => n_285, A2 => n_343, B1 => n_284, B2 => FE_PHN132_framebuffer_buf_28_2316, ZN => n_281);
  g23430 : MOAI22D0BWP7T port map(A1 => n_285, A2 => n_341, B1 => n_284, B2 => FE_PHN128_framebuffer_buf_29_2317, ZN => n_280);
  g23431 : MOAI22D0BWP7T port map(A1 => n_285, A2 => n_339, B1 => n_284, B2 => FE_PHN76_framebuffer_buf_30_2318, ZN => n_279);
  g23434 : MOAI22D0BWP7T port map(A1 => n_285, A2 => n_336, B1 => n_284, B2 => FE_PHN120_framebuffer_buf_31_2319, ZN => n_278);
  g23336 : MOAI22D0BWP7T port map(A1 => n_276, A2 => n_353, B1 => n_275, B2 => framebuffer_buf_128_2416, ZN => n_277);
  g23337 : MOAI22D0BWP7T port map(A1 => n_276, A2 => n_350, B1 => n_275, B2 => FE_PHN164_framebuffer_buf_129_2417, ZN => n_274);
  g23338 : MOAI22D0BWP7T port map(A1 => n_276, A2 => n_347, B1 => n_275, B2 => framebuffer_buf_130_2418, ZN => n_273);
  g23440 : MOAI22D0BWP7T port map(A1 => n_271, A2 => n_353, B1 => n_270, B2 => FE_PHN7_framebuffer_buf_152_2440, ZN => n_272);
  g23339 : MOAI22D0BWP7T port map(A1 => n_276, A2 => n_345, B1 => n_275, B2 => FE_PHN170_framebuffer_buf_131_2419, ZN => n_269);
  g23441 : MOAI22D0BWP7T port map(A1 => n_271, A2 => n_350, B1 => n_270, B2 => FE_PHN185_framebuffer_buf_153_2441, ZN => n_268);
  g23442 : MOAI22D0BWP7T port map(A1 => n_271, A2 => n_347, B1 => n_270, B2 => FE_PHN118_framebuffer_buf_154_2442, ZN => n_267);
  g23443 : MOAI22D0BWP7T port map(A1 => n_271, A2 => n_343, B1 => n_270, B2 => FE_PHN97_framebuffer_buf_156_2444, ZN => n_266);
  g23340 : MOAI22D0BWP7T port map(A1 => n_276, A2 => n_343, B1 => n_275, B2 => FE_PHN91_framebuffer_buf_132_2420, ZN => n_265);
  g23444 : MOAI22D0BWP7T port map(A1 => n_271, A2 => n_341, B1 => n_270, B2 => FE_PHN44_framebuffer_buf_157_2445, ZN => n_264);
  g23445 : MOAI22D0BWP7T port map(A1 => n_262, A2 => n_353, B1 => n_261, B2 => FE_PHN64_framebuffer_buf_64_2352, ZN => n_263);
  g23446 : MOAI22D0BWP7T port map(A1 => n_262, A2 => n_350, B1 => n_261, B2 => FE_PHN16_framebuffer_buf_65_2353, ZN => n_260);
  g23447 : MOAI22D0BWP7T port map(A1 => n_262, A2 => n_347, B1 => n_261, B2 => FE_PHN183_framebuffer_buf_66_2354, ZN => n_259);
  g23342 : MOAI22D0BWP7T port map(A1 => n_251, A2 => n_353, B1 => n_250, B2 => FE_PHN38_framebuffer_buf_144_2432, ZN => n_258);
  g23448 : MOAI22D0BWP7T port map(A1 => n_262, A2 => n_345, B1 => n_261, B2 => FE_PHN12_framebuffer_buf_67_2355, ZN => n_257);
  g23341 : MOAI22D0BWP7T port map(A1 => n_276, A2 => n_341, B1 => n_275, B2 => FE_PHN6_framebuffer_buf_133_2421, ZN => n_256);
  g23449 : MOAI22D0BWP7T port map(A1 => n_318, A2 => n_341, B1 => n_317, B2 => FE_PHN43_framebuffer_buf_53_2341, ZN => n_255);
  g23451 : MOAI22D0BWP7T port map(A1 => n_262, A2 => n_339, B1 => n_261, B2 => FE_PHN84_framebuffer_buf_70_2358, ZN => n_254);
  g23450 : MOAI22D0BWP7T port map(A1 => n_262, A2 => n_341, B1 => n_261, B2 => FE_PHN53_framebuffer_buf_69_2357, ZN => n_253);
  g23343 : MOAI22D0BWP7T port map(A1 => n_251, A2 => n_350, B1 => n_250, B2 => FE_PHN105_framebuffer_buf_145_2433, ZN => n_252);
  g23381 : MOAI22D0BWP7T port map(A1 => n_337, A2 => n_341, B1 => n_335, B2 => FE_PHN65_framebuffer_buf_125_2413, ZN => n_249);
  g23452 : MOAI22D0BWP7T port map(A1 => n_262, A2 => n_336, B1 => n_261, B2 => FE_PHN136_framebuffer_buf_71_2359, ZN => n_248);
  g23453 : MOAI22D0BWP7T port map(A1 => n_246, A2 => n_353, B1 => n_245, B2 => FE_PHN48_framebuffer_buf_72_2360, ZN => n_247);
  g23345 : MOAI22D0BWP7T port map(A1 => n_251, A2 => n_345, B1 => n_250, B2 => FE_PHN2_framebuffer_buf_147_2435, ZN => n_244);
  g23454 : MOAI22D0BWP7T port map(A1 => n_246, A2 => n_350, B1 => n_245, B2 => FE_PHN124_framebuffer_buf_73_2361, ZN => n_243);
  g23346 : MOAI22D0BWP7T port map(A1 => n_251, A2 => n_343, B1 => n_250, B2 => FE_PHN13_framebuffer_buf_148_2436, ZN => n_242);
  g23455 : MOAI22D0BWP7T port map(A1 => n_246, A2 => n_347, B1 => n_245, B2 => FE_PHN17_framebuffer_buf_74_2362, ZN => n_241);
  g23456 : MOAI22D0BWP7T port map(A1 => n_230, A2 => n_353, B1 => n_229, B2 => FE_PHN60_framebuffer_buf_0_2288, ZN => n_240);
  g23457 : MOAI22D0BWP7T port map(A1 => n_246, A2 => n_345, B1 => n_245, B2 => FE_PHN151_framebuffer_buf_75_2363, ZN => n_239);
  g23347 : MOAI22D0BWP7T port map(A1 => n_251, A2 => n_341, B1 => n_250, B2 => FE_PHN21_framebuffer_buf_149_2437, ZN => n_238);
  g23458 : MOAI22D0BWP7T port map(A1 => n_246, A2 => n_343, B1 => n_245, B2 => FE_PHN81_framebuffer_buf_76_2364, ZN => n_237);
  g23459 : MOAI22D0BWP7T port map(A1 => n_246, A2 => n_341, B1 => n_245, B2 => FE_PHN15_framebuffer_buf_77_2365, ZN => n_236);
  g23461 : MOAI22D0BWP7T port map(A1 => n_246, A2 => n_336, B1 => n_245, B2 => FE_PHN20_framebuffer_buf_79_2367, ZN => n_235);
  g23349 : MOAI22D0BWP7T port map(A1 => n_233, A2 => n_350, B1 => n_232, B2 => FE_PHN66_framebuffer_buf_41_2329, ZN => n_234);
  g23463 : MOAI22D0BWP7T port map(A1 => n_230, A2 => n_350, B1 => n_229, B2 => FE_PHN166_framebuffer_buf_1_2289, ZN => n_231);
  g23350 : MOAI22D0BWP7T port map(A1 => n_233, A2 => n_347, B1 => n_232, B2 => FE_PHN140_framebuffer_buf_42_2330, ZN => n_228);
  g23464 : MOAI22D0BWP7T port map(A1 => n_230, A2 => n_347, B1 => n_229, B2 => FE_PHN69_framebuffer_buf_2_2290, ZN => n_227);
  g23465 : MOAI22D0BWP7T port map(A1 => n_225, A2 => n_350, B1 => n_224, B2 => FE_PHN102_framebuffer_buf_81_2369, ZN => n_226);
  g23466 : MOAI22D0BWP7T port map(A1 => n_225, A2 => n_347, B1 => n_224, B2 => framebuffer_buf_82_2370, ZN => n_223);
  g23467 : MOAI22D0BWP7T port map(A1 => n_230, A2 => n_345, B1 => n_229, B2 => framebuffer_buf_3_2291, ZN => n_222);
  g23351 : MOAI22D0BWP7T port map(A1 => n_233, A2 => n_343, B1 => n_232, B2 => framebuffer_buf_44_2332, ZN => n_221);
  g23352 : MOAI22D0BWP7T port map(A1 => n_233, A2 => n_341, B1 => n_232, B2 => FE_PHN90_framebuffer_buf_45_2333, ZN => n_220);
  g23468 : MOAI22D0BWP7T port map(A1 => n_225, A2 => n_345, B1 => n_224, B2 => FE_PHN10_framebuffer_buf_83_2371, ZN => n_219);
  g23353 : MOAI22D0BWP7T port map(A1 => n_213, A2 => n_353, B1 => n_212, B2 => FE_PHN168_framebuffer_buf_56_2344, ZN => n_218);
  g23469 : MOAI22D0BWP7T port map(A1 => n_225, A2 => n_343, B1 => n_224, B2 => FE_PHN145_framebuffer_buf_84_2372, ZN => n_217);
  g23470 : MOAI22D0BWP7T port map(A1 => n_230, A2 => n_343, B1 => n_229, B2 => framebuffer_buf_4_2292, ZN => n_216);
  g23471 : MOAI22D0BWP7T port map(A1 => n_225, A2 => n_341, B1 => n_224, B2 => FE_PHN114_framebuffer_buf_85_2373, ZN => n_215);
  g23354 : MOAI22D0BWP7T port map(A1 => n_213, A2 => n_350, B1 => n_212, B2 => FE_PHN11_framebuffer_buf_57_2345, ZN => n_214);
  g23472 : MOAI22D0BWP7T port map(A1 => n_225, A2 => n_339, B1 => n_224, B2 => FE_PHN100_framebuffer_buf_86_2374, ZN => n_211);
  g23473 : MOAI22D0BWP7T port map(A1 => n_225, A2 => n_336, B1 => n_224, B2 => FE_PHN72_framebuffer_buf_87_2375, ZN => n_210);
  g23474 : MOAI22D0BWP7T port map(A1 => n_206, A2 => n_353, B1 => n_205, B2 => FE_PHN89_framebuffer_buf_88_2376, ZN => n_209);
  g23355 : MOAI22D0BWP7T port map(A1 => n_213, A2 => n_347, B1 => n_212, B2 => FE_PHN57_framebuffer_buf_58_2346, ZN => n_208);
  g23475 : MOAI22D0BWP7T port map(A1 => n_206, A2 => n_350, B1 => n_205, B2 => FE_PHN31_framebuffer_buf_89_2377, ZN => n_207);
  g23356 : MOAI22D0BWP7T port map(A1 => n_213, A2 => n_345, B1 => n_212, B2 => framebuffer_buf_59_2347, ZN => n_204);
  g23476 : MOAI22D0BWP7T port map(A1 => n_230, A2 => n_341, B1 => n_229, B2 => FE_PHN101_framebuffer_buf_5_2293, ZN => n_203);
  g23477 : MOAI22D0BWP7T port map(A1 => n_230, A2 => n_339, B1 => n_229, B2 => FE_PHN67_framebuffer_buf_6_2294, ZN => n_202);
  g23357 : MOAI22D0BWP7T port map(A1 => n_213, A2 => n_343, B1 => n_212, B2 => FE_PHN138_framebuffer_buf_60_2348, ZN => n_201);
  g23478 : MOAI22D0BWP7T port map(A1 => n_206, A2 => n_347, B1 => n_205, B2 => FE_PHN9_framebuffer_buf_90_2378, ZN => n_200);
  g23479 : MOAI22D0BWP7T port map(A1 => n_206, A2 => n_345, B1 => n_205, B2 => FE_PHN79_framebuffer_buf_91_2379, ZN => n_199);
  g23358 : MOAI22D0BWP7T port map(A1 => n_213, A2 => n_341, B1 => n_212, B2 => FE_PHN40_framebuffer_buf_61_2349, ZN => n_198);
  g23480 : MOAI22D0BWP7T port map(A1 => n_230, A2 => n_336, B1 => n_229, B2 => FE_PHN92_framebuffer_buf_7_2295, ZN => n_197);
  g23481 : MOAI22D0BWP7T port map(A1 => n_206, A2 => n_343, B1 => n_205, B2 => FE_PHN182_framebuffer_buf_92_2380, ZN => n_196);
  g23482 : MOAI22D0BWP7T port map(A1 => n_206, A2 => n_341, B1 => n_205, B2 => FE_PHN163_framebuffer_buf_93_2381, ZN => n_195);
  g23360 : MOAI22D0BWP7T port map(A1 => n_276, A2 => n_339, B1 => n_275, B2 => FE_PHN172_framebuffer_buf_134_2422, ZN => n_194);
  g23483 : MOAI22D0BWP7T port map(A1 => n_206, A2 => n_339, B1 => n_205, B2 => FE_PHN62_framebuffer_buf_94_2382, ZN => n_193);
  g23484 : MOAI22D0BWP7T port map(A1 => n_206, A2 => n_336, B1 => n_205, B2 => FE_PHN63_framebuffer_buf_95_2383, ZN => n_192);
  g23359 : MOAI22D0BWP7T port map(A1 => n_233, A2 => n_345, B1 => n_232, B2 => FE_PHN152_framebuffer_buf_43_2331, ZN => n_191);
  g23485 : MOAI22D0BWP7T port map(A1 => n_187, A2 => n_353, B1 => n_186, B2 => FE_PHN54_framebuffer_buf_96_2384, ZN => n_190);
  g23361 : MOAI22D0BWP7T port map(A1 => n_318, A2 => n_347, B1 => n_317, B2 => FE_PHN165_framebuffer_buf_50_2338, ZN => n_189);
  g23486 : MOAI22D0BWP7T port map(A1 => n_187, A2 => n_350, B1 => n_186, B2 => FE_PHN46_framebuffer_buf_97_2385, ZN => n_188);
  g23362 : MOAI22D0BWP7T port map(A1 => n_251, A2 => n_339, B1 => n_250, B2 => framebuffer_buf_150_2438, ZN => n_185);
  g23487 : MOAI22D0BWP7T port map(A1 => n_187, A2 => n_347, B1 => n_186, B2 => framebuffer_buf_98_2386, ZN => n_184);
  g23488 : MOAI22D0BWP7T port map(A1 => n_187, A2 => n_345, B1 => n_186, B2 => framebuffer_buf_99_2387, ZN => n_183);
  g23489 : MOAI22D0BWP7T port map(A1 => n_187, A2 => n_343, B1 => n_186, B2 => FE_PHN70_framebuffer_buf_100_2388, ZN => n_182);
  g23363 : MOAI22D0BWP7T port map(A1 => n_251, A2 => n_336, B1 => n_250, B2 => FE_PHN177_framebuffer_buf_151_2439, ZN => n_181);
  g23490 : MOAI22D0BWP7T port map(A1 => n_187, A2 => n_341, B1 => n_186, B2 => FE_PHN55_framebuffer_buf_101_2389, ZN => n_180);
  g23491 : MOAI22D0BWP7T port map(A1 => n_187, A2 => n_339, B1 => n_186, B2 => FE_PHN117_framebuffer_buf_102_2390, ZN => n_179);
  g23492 : MOAI22D0BWP7T port map(A1 => n_187, A2 => n_336, B1 => n_186, B2 => FE_PHN56_framebuffer_buf_103_2391, ZN => n_178);
  g23493 : MOAI22D0BWP7T port map(A1 => n_301, A2 => n_353, B1 => n_300, B2 => FE_PHN131_framebuffer_buf_16_2304, ZN => n_177);
  g23364 : MOAI22D0BWP7T port map(A1 => n_233, A2 => n_339, B1 => n_232, B2 => FE_PHN109_framebuffer_buf_46_2334, ZN => n_176);
  g23365 : MOAI22D0BWP7T port map(A1 => n_233, A2 => n_336, B1 => n_232, B2 => framebuffer_buf_47_2335, ZN => n_175);
  g23366 : MOAI22D0BWP7T port map(A1 => n_213, A2 => n_339, B1 => n_212, B2 => FE_PHN142_framebuffer_buf_62_2350, ZN => n_174);
  g23367 : MOAI22D0BWP7T port map(A1 => n_213, A2 => n_336, B1 => n_212, B2 => FE_PHN78_framebuffer_buf_63_2351, ZN => n_173);
  g23368 : MOAI22D0BWP7T port map(A1 => n_170, A2 => n_353, B1 => n_169, B2 => FE_PHN157_framebuffer_buf_104_2392, ZN => n_172);
  g23369 : MOAI22D0BWP7T port map(A1 => n_170, A2 => n_350, B1 => n_169, B2 => FE_PHN180_framebuffer_buf_105_2393, ZN => n_171);
  g23370 : MOAI22D0BWP7T port map(A1 => n_170, A2 => n_347, B1 => n_169, B2 => FE_PHN47_framebuffer_buf_106_2394, ZN => n_168);
  g23371 : MOAI22D0BWP7T port map(A1 => n_170, A2 => n_345, B1 => n_169, B2 => FE_PHN146_framebuffer_buf_107_2395, ZN => n_167);
  g23372 : MOAI22D0BWP7T port map(A1 => n_170, A2 => n_343, B1 => n_169, B2 => FE_PHN153_framebuffer_buf_108_2396, ZN => n_166);
  g23373 : MOAI22D0BWP7T port map(A1 => n_170, A2 => n_341, B1 => n_169, B2 => framebuffer_buf_109_2397, ZN => n_165);
  g23374 : MOAI22D0BWP7T port map(A1 => n_170, A2 => n_336, B1 => n_169, B2 => FE_PHN71_framebuffer_buf_111_2399, ZN => n_164);
  g23375 : MOAI22D0BWP7T port map(A1 => n_170, A2 => n_339, B1 => n_169, B2 => FE_PHN52_framebuffer_buf_110_2398, ZN => n_163);
  g23376 : MOAI22D0BWP7T port map(A1 => n_337, A2 => n_353, B1 => n_335, B2 => FE_PHN75_framebuffer_buf_120_2408, ZN => n_162);
  g23377 : MOAI22D0BWP7T port map(A1 => n_337, A2 => n_350, B1 => n_335, B2 => FE_PHN29_framebuffer_buf_121_2409, ZN => n_161);
  g23378 : MOAI22D0BWP7T port map(A1 => n_337, A2 => n_347, B1 => n_335, B2 => FE_PHN45_framebuffer_buf_122_2410, ZN => n_160);
  g23379 : MOAI22D0BWP7T port map(A1 => n_337, A2 => n_345, B1 => n_335, B2 => FE_PHN179_framebuffer_buf_123_2411, ZN => n_159);
  g23380 : MOAI22D0BWP7T port map(A1 => n_337, A2 => n_343, B1 => n_335, B2 => FE_PHN96_framebuffer_buf_124_2412, ZN => n_158);
  g23344 : MOAI22D0BWP7T port map(A1 => n_251, A2 => n_347, B1 => n_250, B2 => FE_PHN80_framebuffer_buf_146_2434, ZN => n_157);
  new_counter_reg_5 : LHQD1BWP7T port map(D => n_146, E => n_396, Q => new_counter(5));
  g23109 : OAI21D0BWP7T port map(A1 => n_150, A2 => counter(6), B => n_148, ZN => n_156);
  state_reg_1 : DFKCNQD1BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_135, Q => state(1));
  g23110 : ND2D0BWP7T port map(A1 => n_147, A2 => counter(6), ZN => n_155);
  state_reg_0 : DFKCNQD1BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_123, Q => state(0));
  counter_reg_3 : DFKCNQD1BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => new_counter(3), Q => counter(3));
  g23515 : OAI211D1BWP7T port map(A1 => n_154, A2 => n_139, B => n_153, C => n_152, ZN => n_385);
  g23514 : OAI211D1BWP7T port map(A1 => n_154, A2 => n_141, B => n_153, C => n_152, ZN => n_377);
  g23498 : OAI211D0BWP7T port map(A1 => n_154, A2 => n_140, B => n_153, C => n_149, ZN => n_391);
  g23532 : OAI21D0BWP7T port map(A1 => n_129, A2 => n_143, B => n_142, ZN => n_366);
  g23497 : OAI211D0BWP7T port map(A1 => sqi_finished, A2 => n_150, B => n_149, C => n_57, ZN => n_151);
  new_counter_reg_4 : LHQD1BWP7T port map(D => n_120, E => n_396, Q => new_counter(4));
  g23115 : INVD0BWP7T port map(I => n_147, ZN => n_148);
  g23108 : OAI22D0BWP7T port map(A1 => n_136, A2 => n_145, B1 => n_144, B2 => counter(5), ZN => n_146);
  g23525 : OAI21D0BWP7T port map(A1 => n_127, A2 => n_143, B => n_142, ZN => n_270);
  g23516 : OAI21D0BWP7T port map(A1 => n_118, A2 => n_143, B => n_142, ZN => n_275);
  counter_reg_1 : DFKCNQD1BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => new_counter(1), Q => counter(1));
  g23517 : OAI21D0BWP7T port map(A1 => n_126, A2 => n_143, B => n_142, ZN => n_250);
  g23518 : OAI21D0BWP7T port map(A1 => n_86, A2 => n_143, B => n_142, ZN => n_232);
  g23519 : OAI21D0BWP7T port map(A1 => n_90, A2 => n_143, B => n_142, ZN => n_212);
  g23521 : OAI21D0BWP7T port map(A1 => n_89, A2 => n_143, B => n_142, ZN => n_169);
  counter_reg_2 : DFKCNQD1BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => new_counter(2), Q => counter(2));
  g23526 : OAI21D0BWP7T port map(A1 => n_97, A2 => n_143, B => n_142, ZN => n_284);
  g23527 : OAI21D0BWP7T port map(A1 => n_100, A2 => n_143, B => n_142, ZN => n_303);
  g23528 : OAI21D0BWP7T port map(A1 => n_101, A2 => n_143, B => n_142, ZN => n_224);
  g23529 : OAI21D0BWP7T port map(A1 => n_85, A2 => n_143, B => n_142, ZN => n_261);
  g23530 : OAI21D0BWP7T port map(A1 => n_87, A2 => n_143, B => n_142, ZN => n_186);
  g23531 : OAI21D0BWP7T port map(A1 => n_78, A2 => n_143, B => n_142, ZN => n_335);
  g23533 : OAI21D0BWP7T port map(A1 => n_77, A2 => n_143, B => n_142, ZN => n_245);
  g23534 : OAI21D0BWP7T port map(A1 => n_141, A2 => n_143, B => n_142, ZN => n_300);
  g23535 : OAI21D0BWP7T port map(A1 => n_96, A2 => n_143, B => n_142, ZN => n_205);
  g23536 : OAI21D0BWP7T port map(A1 => n_140, A2 => n_143, B => n_142, ZN => n_229);
  g23537 : OAI21D0BWP7T port map(A1 => n_139, A2 => n_143, B => n_142, ZN => n_349);
  g23538 : OAI21D0BWP7T port map(A1 => n_93, A2 => n_143, B => n_142, ZN => n_329);
  g23539 : OAI21D0BWP7T port map(A1 => n_88, A2 => n_143, B => n_142, ZN => n_317);
  g23500 : INVD5BWP7T port map(I => n_407, ZN => sqi_data_out(2));
  g23502 : INVD5BWP7T port map(I => n_406, ZN => sqi_data_out(1));
  g23116 : OAI21D0BWP7T port map(A1 => n_150, A2 => counter(5), B => n_136, ZN => n_147);
  state_reg_3 : DFQD1BWP7T port map(CP => CTS_13, D => n_117, Q => state(3));
  g23508 : ND2D0BWP7T port map(A1 => n_116, A2 => n_98, ZN => n_135);
  g23506 : INVD5BWP7T port map(I => n_404, ZN => sqi_data_out(5));
  g23504 : INVD5BWP7T port map(I => n_405, ZN => sqi_data_out(3));
  g23512 : INVD5BWP7T port map(I => n_403, ZN => sqi_data_out(4));
  g23520 : IND4D0BWP7T port map(A1 => n_128, B1 => n_52, B2 => n_92, B3 => n_150, ZN => n_397);
  new_counter_reg_3 : LHQD1BWP7T port map(D => n_104, E => n_396, Q => new_counter(3));
  g23553 : INVD5BWP7T port map(I => n_401, ZN => sqi_data_out(6));
  g23555 : INVD5BWP7T port map(I => n_400, ZN => sqi_data_out(7));
  g23563 : INVD0BWP7T port map(I => n_1522, ZN => n_129);
  g23556 : NR2XD0BWP7T port map(A1 => n_128, A2 => n_29, ZN => n_153);
  g23560 : INVD1BWP7T port map(I => n_127, ZN => n_271);
  g23562 : INVD1BWP7T port map(I => n_126, ZN => n_251);
  g23582 : NR2XD0BWP7T port map(A1 => n_301, A2 => n_154, ZN => n_376);
  g23551 : NR3D1BWP7T port map(A1 => n_128, A2 => n_33, A3 => n_121, ZN => n_142);
  g23541 : INVD5BWP7T port map(I => n_402, ZN => sqi_data_out(0));
  sqi_data_out_reg_2 : LHD1BWP7T port map(D => n_110, E => n_124, Q => UNCONNECTED, QN => n_407);
  sqi_data_out_reg_1 : LHD1BWP7T port map(D => n_109, E => n_124, Q => UNCONNECTED0, QN => n_406);
  sqi_data_out_reg_3 : LHD1BWP7T port map(D => n_103, E => n_124, Q => UNCONNECTED1, QN => n_405);
  sqi_data_out_reg_5 : LHD1BWP7T port map(D => n_105, E => n_124, Q => UNCONNECTED2, QN => n_404);
  g23509 : IND4D0BWP7T port map(A1 => n_115, B1 => n_35, B2 => n_47, B3 => n_95, ZN => n_123);
  sqi_data_out_reg_4 : LHD1BWP7T port map(D => n_106, E => n_124, Q => UNCONNECTED3, QN => n_403);
  g23523 : AOI22D0BWP7T port map(A1 => n_113, A2 => n_121, B1 => n_80, B2 => sqi_finished, ZN => n_122);
  g23117 : OAI22D0BWP7T port map(A1 => n_112, A2 => n_45, B1 => n_81, B2 => n_111, ZN => n_120);
  state_reg_2 : DFQD1BWP7T port map(CP => CTS_13, D => n_102, Q => state(2));
  sqi_data_out_reg_7 : LHD1BWP7T port map(D => n_43, E => n_124, Q => UNCONNECTED4, QN => n_400);
  sqi_data_out_reg_6 : LHD1BWP7T port map(D => n_67, E => n_124, Q => UNCONNECTED5, QN => n_401);
  g23572 : NR2XD0BWP7T port map(A1 => n_119, A2 => counter(0), ZN => n_126);
  g23570 : NR2XD0BWP7T port map(A1 => n_119, A2 => n_22, ZN => n_127);
  g23561 : INVD1BWP7T port map(I => n_118, ZN => n_276);
  g23583 : NR2D0BWP7T port map(A1 => n_230, A2 => n_154, ZN => n_390);
  g23510 : OR4D1BWP7T port map(A1 => reset, A2 => n_5, A3 => n_114, A4 => n_75, Z => n_117);
  new_counter_reg_2 : LHQD1BWP7T port map(D => n_63, E => n_396, Q => new_counter(2));
  new_counter_reg_1 : LHQD1BWP7T port map(D => n_74, E => n_396, Q => new_counter(1));
  g23542 : NR4D0BWP7T port map(A1 => n_115, A2 => n_65, A3 => n_114, A4 => n_46, ZN => n_116);
  sqi_data_out_reg_0 : LHD1BWP7T port map(D => n_94, E => n_124, Q => UNCONNECTED6, QN => n_402);
  g23543 : IND2D0BWP7T port map(A1 => n_113, B1 => n_121, ZN => n_149);
  g23301 : AN2D1BWP7T port map(A1 => n_112, A2 => n_111, Z => n_136);
  g23584 : NR2XD0BWP7T port map(A1 => n_351, A2 => n_154, ZN => n_384);
  g23547 : AO22D0BWP7T port map(A1 => n_108, A2 => row_buf(2), B1 => calc_buf_in(1), B2 => n_107, Z => n_110);
  g23548 : AO22D0BWP7T port map(A1 => n_108, A2 => row_buf(1), B1 => calc_buf_in(0), B2 => n_107, Z => n_109);
  g23549 : AO22D0BWP7T port map(A1 => n_108, A2 => row_buf(4), B1 => calc_buf_in(3), B2 => n_107, Z => n_106);
  g23550 : AO22D0BWP7T port map(A1 => n_108, A2 => row_buf(5), B1 => calc_buf_in(4), B2 => n_107, Z => n_105);
  g23310 : MOAI22D0BWP7T port map(A1 => n_55, A2 => n_150, B1 => n_79, B2 => counter(3), ZN => n_104);
  g23546 : AO22D0BWP7T port map(A1 => n_108, A2 => row_buf(3), B1 => calc_buf_in(2), B2 => n_107, Z => n_103);
  g23571 : NR2XD0BWP7T port map(A1 => n_83, A2 => counter(0), ZN => n_118);
  g23513 : ND4D0BWP7T port map(A1 => n_91, A2 => n_51, A3 => n_143, A4 => FE_OFN0_FE_DBTN0_reset, ZN => n_102);
  g23587 : INVD0BWP7T port map(I => n_225, ZN => n_101);
  g23588 : INVD0BWP7T port map(I => n_1523, ZN => n_100);
  g23211 : NR2D0BWP7T port map(A1 => n_144, A2 => counter(7), ZN => n_99);
  g23580 : ND2D1BWP7T port map(A1 => n_66, A2 => n_98, ZN => n_128);
  g23609 : INVD1BWP7T port map(I => n_97, ZN => n_285);
  g23610 : INVD1BWP7T port map(I => n_96, ZN => n_206);
  g23612 : INVD1BWP7T port map(I => n_141, ZN => n_301);
  g23577 : AOI31D0BWP7T port map(A1 => n_40, A2 => state(1), A3 => sqi_finished, B => n_50, ZN => n_95);
  g23557 : INR2D0BWP7T port map(A1 => row_buf(0), B1 => n_98, ZN => n_94);
  g23595 : ND2D1BWP7T port map(A1 => n_82, A2 => n_61, ZN => n_119);
  g23558 : NR3D0BWP7T port map(A1 => n_59, A2 => counter(1), A3 => counter(2), ZN => n_113);
  g23581 : ND2D0BWP7T port map(A1 => n_58, A2 => n_98, ZN => n_124);
  g23585 : INVD1BWP7T port map(I => n_93, ZN => n_330);
  g23545 : OAI211D0BWP7T port map(A1 => n_152, A2 => n_92, B => n_91, C => n_150, ZN => n_396);
  g23590 : INVD1BWP7T port map(I => n_90, ZN => n_213);
  g23591 : INVD1BWP7T port map(I => n_89, ZN => n_170);
  g23593 : INVD1BWP7T port map(I => n_88, ZN => n_318);
  g23594 : INVD1BWP7T port map(I => n_87, ZN => n_187);
  g23589 : INVD1BWP7T port map(I => n_86, ZN => n_233);
  g23586 : INVD0BWP7T port map(I => n_262, ZN => n_85);
  g23622 : INR2XD0BWP7T port map(A1 => n_82, B1 => n_70, ZN => n_97);
  g23623 : INR2XD0BWP7T port map(A1 => n_82, B1 => n_68, ZN => n_96);
  g23307 : AOI21D0BWP7T port map(A1 => n_81, A2 => n_80, B => n_79, ZN => n_112);
  g23625 : INR2XD0BWP7T port map(A1 => n_82, B1 => n_72, ZN => n_141);
  g23592 : INVD1BWP7T port map(I => n_78, ZN => n_337);
  g23611 : INVD1BWP7T port map(I => n_77, ZN => n_246);
  g23614 : INVD1BWP7T port map(I => n_139, ZN => n_351);
  g23613 : INVD1BWP7T port map(I => n_140, ZN => n_230);
  g23600 : ND2D1BWP7T port map(A1 => n_82, A2 => n_76, ZN => n_225);
  g23574 : OAI211D1BWP7T port map(A1 => n_12, A2 => n_9, B => n_73, C => n_6, ZN => n_75);
  g23576 : MOAI22D0BWP7T port map(A1 => n_150, A2 => n_17, B1 => n_79, B2 => counter(1), ZN => n_74);
  g23559 : OAI211D1BWP7T port map(A1 => ce, A2 => n_64, B => n_73, C => n_32, ZN => n_115);
  g23598 : NR2D1BWP7T port map(A1 => n_71, A2 => n_72, ZN => n_93);
  g23606 : NR2D1BWP7T port map(A1 => n_69, A2 => n_72, ZN => n_88);
  g23602 : NR2D1BWP7T port map(A1 => n_71, A2 => n_70, ZN => n_86);
  g23603 : NR2D1BWP7T port map(A1 => n_69, A2 => n_70, ZN => n_90);
  g23604 : NR2XD0BWP7T port map(A1 => n_71, A2 => n_68, ZN => n_89);
  g23605 : NR2XD0BWP7T port map(A1 => n_69, A2 => n_68, ZN => n_78);
  g23599 : ND2D1BWP7T port map(A1 => n_62, A2 => n_76, ZN => n_262);
  g23620 : AO22D0BWP7T port map(A1 => n_107, A2 => calc_buf_in(5), B1 => calc_buf_in(0), B2 => n_108, Z => n_67);
  g23617 : AOI211XD0BWP7T port map(A1 => n_10, A2 => state(1), B => n_34, C => n_107, ZN => n_66);
  g23616 : OAI211D1BWP7T port map(A1 => mode, A2 => n_64, B => n_51, C => n_42, ZN => n_65);
  g23522 : MOAI22D0BWP7T port map(A1 => n_39, A2 => n_150, B1 => n_79, B2 => counter(2), ZN => n_63);
  g23621 : ND2D1BWP7T port map(A1 => n_62, A2 => n_61, ZN => n_83);
  g23624 : INR2XD0BWP7T port map(A1 => n_62, B1 => n_68, ZN => n_77);
  g23607 : INR2XD0BWP7T port map(A1 => n_76, B1 => n_71, ZN => n_87);
  g23627 : INR2XD0BWP7T port map(A1 => n_62, B1 => n_70, ZN => n_139);
  g23308 : IND3D0BWP7T port map(A1 => n_81, B1 => counter(4), B2 => n_80, ZN => n_144);
  g23626 : INR2XD0BWP7T port map(A1 => n_62, B1 => n_72, ZN => n_140);
  row_buf_reg_1 : DFKCNQD1BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => new_row_buf(1), Q => row_buf(1));
  row_buf_reg_2 : DFKCNQD1BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => new_row_buf(2), Q => row_buf(2));
  row_buf_reg_0 : DFKCNQD1BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => new_row_buf(0), Q => row_buf(0));
  g23618 : IND4D0BWP7T port map(A1 => n_72, B1 => n_7, B2 => n_4, B3 => n_20, ZN => n_59);
  g23619 : OAI21D0BWP7T port map(A1 => n_15, A2 => n_56, B => n_107, ZN => n_58);
  g23579 : OAI222D0BWP7T port map(A1 => n_48, A2 => n_57, B1 => n_56, B2 => n_49, C1 => n_41, C2 => n_25, ZN => n_114);
  g23524 : MAOI22D0BWP7T port map(A1 => n_54, A2 => counter(3), B1 => n_54, B2 => counter(3), ZN => n_55);
  row_buf_reg_3 : DFKCNQD1BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => new_row_buf(3), Q => row_buf(3));
  row_buf_reg_4 : DFKCNQD1BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => new_row_buf(4), Q => row_buf(4));
  row_buf_reg_5 : DFKCNQD1BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => new_row_buf(5), Q => row_buf(5));
  g23615 : OAI22D0BWP7T port map(A1 => n_49, A2 => n_26, B1 => n_143, B2 => sqi_finished, ZN => n_50);
  g23646 : NR2XD0BWP7T port map(A1 => n_37, A2 => counter(2), ZN => n_82);
  g23578 : AOI22D0BWP7T port map(A1 => n_48, A2 => n_21, B1 => n_18, B2 => ce, ZN => n_91);
  g23544 : IND2D0BWP7T port map(A1 => n_54, B1 => counter(3), ZN => n_81);
  g23635 : INR2XD0BWP7T port map(A1 => n_44, B1 => counter(2), ZN => n_62);
  g23636 : INVD0BWP7T port map(I => n_46, ZN => n_47);
  g23641 : ND2D0BWP7T port map(A1 => n_80, A2 => n_45, ZN => n_111);
  g23644 : ND2D1BWP7T port map(A1 => n_44, A2 => counter(2), ZN => n_71);
  g23645 : ND2D1BWP7T port map(A1 => n_36, A2 => counter(2), ZN => n_69);
  g23634 : INR2D0BWP7T port map(A1 => calc_buf_in(1), B1 => n_98, ZN => n_43);
  g23638 : AOI22D0BWP7T port map(A1 => n_11, A2 => n_41, B1 => n_13, B2 => n_40, ZN => n_42);
  g23575 : MAOI22D0BWP7T port map(A1 => n_38, A2 => counter(2), B1 => n_38, B2 => counter(2), ZN => n_39);
  g23640 : OAI22D0BWP7T port map(A1 => n_27, A2 => rw, B1 => n_52, B2 => reset, ZN => n_46);
  g23596 : ND2D1BWP7T port map(A1 => n_92, A2 => n_121, ZN => n_73);
  g23647 : INVD0BWP7T port map(I => n_36, ZN => n_37);
  g23660 : INVD0BWP7T port map(I => n_34, ZN => n_35);
  g23666 : ND2D1BWP7T port map(A1 => n_33, A2 => sqi_finished, ZN => n_51);
  g23669 : ND2D0BWP7T port map(A1 => n_57, A2 => n_152, ZN => n_79);
  g23663 : INVD0BWP7T port map(I => n_80, ZN => n_150);
  g23652 : ND2D1BWP7T port map(A1 => n_32, A2 => n_49, ZN => n_107);
  new_row_buf_reg_2 : LNQD1BWP7T port map(D => sqi_data_in(2), EN => n_31, Q => new_row_buf(2));
  new_row_buf_reg_4 : LNQD1BWP7T port map(D => sqi_data_in(4), EN => n_31, Q => new_row_buf(4));
  new_row_buf_reg_3 : LNQD1BWP7T port map(D => sqi_data_in(3), EN => n_31, Q => new_row_buf(3));
  g23649 : INR2XD0BWP7T port map(A1 => counter(1), B1 => n_24, ZN => n_36);
  g23597 : IND2D0BWP7T port map(A1 => n_38, B1 => counter(2), ZN => n_54);
  g23651 : NR2XD0BWP7T port map(A1 => n_30, A2 => counter(0), ZN => n_76);
  g23650 : IND2D1BWP7T port map(A1 => n_30, B1 => counter(0), ZN => n_68);
  g23653 : ND2D1BWP7T port map(A1 => n_29, A2 => sqi_data_in(6), ZN => n_339);
  g23655 : ND2D1BWP7T port map(A1 => n_29, A2 => sqi_data_in(2), ZN => n_347);
  g23656 : ND2D1BWP7T port map(A1 => n_29, A2 => sqi_data_in(4), ZN => n_343);
  g23657 : ND2D1BWP7T port map(A1 => n_29, A2 => sqi_data_in(5), ZN => n_341);
  g23658 : ND2D1BWP7T port map(A1 => n_29, A2 => sqi_data_in(3), ZN => n_345);
  g23654 : ND2D1BWP7T port map(A1 => n_29, A2 => sqi_data_in(0), ZN => n_353);
  new_row_buf_reg_1 : LNQD1BWP7T port map(D => sqi_data_in(1), EN => n_31, Q => new_row_buf(1));
  g23664 : ND2D5BWP7T port map(A1 => n_27, A2 => n_52, ZN => ready);
  new_row_buf_reg_5 : LNQD1BWP7T port map(D => sqi_data_in(5), EN => n_31, Q => new_row_buf(5));
  new_row_buf_reg_0 : LNQD1BWP7T port map(D => sqi_data_in(0), EN => n_31, Q => new_row_buf(0));
  g23661 : INVD0BWP7T port map(I => n_56, ZN => n_26);
  g23667 : ND2D1BWP7T port map(A1 => n_57, A2 => n_25, ZN => n_34);
  g23648 : NR2XD0BWP7T port map(A1 => n_24, A2 => counter(1), ZN => n_44);
  g23670 : ND2D1BWP7T port map(A1 => n_23, A2 => counter(0), ZN => n_70);
  g23671 : ND2D1BWP7T port map(A1 => n_23, A2 => n_22, ZN => n_72);
  g23674 : ND2D0BWP7T port map(A1 => n_143, A2 => n_154, ZN => n_80);
  g23662 : INVD0BWP7T port map(I => n_98, ZN => n_108);
  g23675 : ND2D1BWP7T port map(A1 => n_29, A2 => sqi_data_in(7), ZN => n_336);
  g23659 : ND2D1BWP7T port map(A1 => n_29, A2 => sqi_data_in(1), ZN => n_350);
  g23678 : INVD0BWP7T port map(I => n_57, ZN => n_21);
  g23642 : OA211D0BWP7T port map(A1 => n_45, A2 => n_19, B => n_20, C => n_0, Z => n_48);
  g23680 : INVD0BWP7T port map(I => n_154, ZN => n_33);
  g23643 : ND4D0BWP7T port map(A1 => n_19, A2 => n_20, A3 => n_14, A4 => n_2, ZN => n_92);
  g23668 : NR4D1BWP7T port map(A1 => n_3, A2 => x(4), A3 => x(0), A4 => x(2), ZN => n_56);
  g23677 : INVD0BWP7T port map(I => n_27, ZN => n_18);
  g23665 : MAOI22D0BWP7T port map(A1 => n_16, A2 => counter(1), B1 => n_16, B2 => counter(1), ZN => n_17);
  g23676 : CKND1BWP7T port map(I => n_15, ZN => n_32);
  g23679 : INVD1BWP7T port map(I => n_121, ZN => n_152);
  g23673 : IND3D1BWP7T port map(A1 => state(2), B1 => state(3), B2 => n_8, ZN => n_98);
  g23684 : INR2XD0BWP7T port map(A1 => n_14, B1 => counter(3), ZN => n_23);
  g23682 : ND2D1BWP7T port map(A1 => n_14, A2 => counter(3), ZN => n_30);
  g23681 : ND2D1BWP7T port map(A1 => n_20, A2 => sqi_finished, ZN => n_24);
  g23685 : NR2D1BWP7T port map(A1 => n_64, A2 => state(1), ZN => n_15);
  g23686 : ND2D1BWP7T port map(A1 => n_13, A2 => state(2), ZN => n_49);
  g23689 : INR2D1BWP7T port map(A1 => state(2), B1 => n_12, ZN => n_121);
  g23672 : IND3D0BWP7T port map(A1 => n_12, B1 => sqi_finished, B2 => state(3), ZN => n_31);
  g23696 : INR2D1BWP7T port map(A1 => n_10, B1 => n_12, ZN => n_11);
  g23692 : IAO21D0BWP7T port map(A1 => state(2), A2 => n_41, B => state(3), ZN => n_9);
  g23683 : ND2D1BWP7T port map(A1 => n_40, A2 => state(0), ZN => n_25);
  g23698 : IND2D0BWP7T port map(A1 => n_16, B1 => counter(1), ZN => n_38);
  g23687 : ND2D1BWP7T port map(A1 => n_13, A2 => state(3), ZN => n_27);
  g23688 : IND2D1BWP7T port map(A1 => n_10, B1 => n_8, ZN => n_57);
  g23690 : CKND2D1BWP7T port map(A1 => n_40, A2 => n_8, ZN => n_154);
  g23691 : INVD1BWP7T port map(I => n_143, ZN => n_29);
  g23693 : NR4D0BWP7T port map(A1 => y(5), A2 => y(4), A3 => y(6), A4 => y(7), ZN => n_7);
  g23694 : IND3D0BWP7T port map(A1 => ce, B1 => state(1), B2 => state(3), ZN => n_6);
  g23706 : INVD0BWP7T port map(I => n_52, ZN => n_5);
  g23695 : NR4D0BWP7T port map(A1 => y(1), A2 => y(0), A3 => y(2), A4 => y(3), ZN => n_4);
  g23697 : NR3D0BWP7T port map(A1 => n_45, A2 => counter(3), A3 => counter(7), ZN => n_61);
  g23699 : IND3D1BWP7T port map(A1 => state(1), B1 => state(2), B2 => state(0), ZN => n_143);
  g23708 : OR2D1BWP7T port map(A1 => x(1), A2 => x(3), Z => n_3);
  g23707 : CKND2D1BWP7T port map(A1 => counter(0), A2 => counter(1), ZN => n_2);
  g23700 : NR2XD0BWP7T port map(A1 => counter(3), A2 => counter(2), ZN => n_19);
  g23703 : NR2XD0BWP7T port map(A1 => counter(4), A2 => counter(7), ZN => n_14);
  g23701 : ND2D0BWP7T port map(A1 => counter(0), A2 => sqi_finished, ZN => n_16);
  g23709 : AN2D1BWP7T port map(A1 => state(0), A2 => state(1), Z => n_13);
  g23705 : IND2D1BWP7T port map(A1 => state(0), B1 => state(1), ZN => n_12);
  g23702 : CKND2D1BWP7T port map(A1 => state(0), A2 => state(3), ZN => n_64);
  g23710 : NR2D1BWP7T port map(A1 => state(0), A2 => state(1), ZN => n_8);
  g23711 : IND2D1BWP7T port map(A1 => state(3), B1 => state(2), ZN => n_10);
  g23704 : NR2XD0BWP7T port map(A1 => counter(5), A2 => counter(6), ZN => n_20);
  g23712 : NR2D1BWP7T port map(A1 => state(3), A2 => state(2), ZN => n_40);
  g23713 : ND2D1BWP7T port map(A1 => state(3), A2 => state(2), ZN => n_52);
  g23717 : INVD0BWP7T port map(I => sqi_finished, ZN => n_41);
  drc_bufs23953 : INVD5BWP7T port map(I => n_430, ZN => framebuffer_buf(0));
  drc_bufs23959 : INVD5BWP7T port map(I => n_436, ZN => framebuffer_buf(157));
  drc_bufs23965 : INVD5BWP7T port map(I => n_442, ZN => framebuffer_buf(156));
  drc_bufs23971 : INVD5BWP7T port map(I => n_448, ZN => framebuffer_buf(7));
  drc_bufs23977 : INVD5BWP7T port map(I => n_454, ZN => framebuffer_buf(154));
  drc_bufs23983 : INVD5BWP7T port map(I => n_460, ZN => framebuffer_buf(153));
  drc_bufs23989 : INVD5BWP7T port map(I => n_466, ZN => framebuffer_buf(152));
  drc_bufs23995 : INVD5BWP7T port map(I => n_472, ZN => framebuffer_buf(8));
  drc_bufs24001 : INVD5BWP7T port map(I => n_478, ZN => framebuffer_buf(150));
  drc_bufs24007 : INVD5BWP7T port map(I => n_484, ZN => framebuffer_buf(149));
  drc_bufs24013 : INVD5BWP7T port map(I => n_490, ZN => framebuffer_buf(148));
  drc_bufs24019 : INVD5BWP7T port map(I => n_496, ZN => framebuffer_buf(147));
  drc_bufs24025 : INVD5BWP7T port map(I => n_502, ZN => framebuffer_buf(146));
  drc_bufs24031 : INVD5BWP7T port map(I => n_508, ZN => framebuffer_buf(145));
  drc_bufs24037 : INVD5BWP7T port map(I => n_514, ZN => framebuffer_buf(144));
  drc_bufs24043 : INVD5BWP7T port map(I => n_520, ZN => framebuffer_buf(9));
  drc_bufs24049 : INVD5BWP7T port map(I => n_526, ZN => framebuffer_buf(142));
  drc_bufs24055 : INVD5BWP7T port map(I => n_532, ZN => framebuffer_buf(141));
  drc_bufs24061 : INVD5BWP7T port map(I => n_538, ZN => framebuffer_buf(140));
  drc_bufs24067 : INVD5BWP7T port map(I => n_544, ZN => framebuffer_buf(39));
  drc_bufs24073 : INVD5BWP7T port map(I => n_550, ZN => framebuffer_buf(138));
  drc_bufs24079 : INVD5BWP7T port map(I => n_556, ZN => framebuffer_buf(40));
  drc_bufs24085 : INVD5BWP7T port map(I => n_562, ZN => framebuffer_buf(136));
  drc_bufs24091 : INVD5BWP7T port map(I => n_568, ZN => framebuffer_buf(103));
  drc_bufs24097 : INVD5BWP7T port map(I => n_574, ZN => framebuffer_buf(134));
  drc_bufs24103 : INVD5BWP7T port map(I => n_580, ZN => framebuffer_buf(133));
  drc_bufs24109 : INVD5BWP7T port map(I => n_586, ZN => framebuffer_buf(132));
  drc_bufs24115 : INVD5BWP7T port map(I => n_592, ZN => framebuffer_buf(131));
  drc_bufs24121 : INVD5BWP7T port map(I => n_598, ZN => framebuffer_buf(130));
  drc_bufs24127 : INVD5BWP7T port map(I => n_604, ZN => framebuffer_buf(129));
  drc_bufs24133 : INVD5BWP7T port map(I => n_610, ZN => framebuffer_buf(128));
  drc_bufs24139 : INVD5BWP7T port map(I => n_616, ZN => framebuffer_buf(104));
  drc_bufs24145 : INVD5BWP7T port map(I => n_622, ZN => framebuffer_buf(126));
  drc_bufs24151 : INVD5BWP7T port map(I => n_628, ZN => framebuffer_buf(125));
  drc_bufs24157 : INVD5BWP7T port map(I => n_634, ZN => framebuffer_buf(124));
  drc_bufs24163 : INVD5BWP7T port map(I => n_640, ZN => framebuffer_buf(105));
  drc_bufs24169 : INVD5BWP7T port map(I => n_646, ZN => framebuffer_buf(122));
  drc_bufs24175 : INVD5BWP7T port map(I => n_652, ZN => framebuffer_buf(121));
  drc_bufs24181 : INVD5BWP7T port map(I => n_658, ZN => framebuffer_buf(120));
  drc_bufs24187 : INVD5BWP7T port map(I => n_664, ZN => framebuffer_buf(106));
  drc_bufs24193 : INVD5BWP7T port map(I => n_670, ZN => framebuffer_buf(118));
  drc_bufs24199 : INVD5BWP7T port map(I => n_676, ZN => framebuffer_buf(117));
  drc_bufs24205 : INVD5BWP7T port map(I => n_682, ZN => framebuffer_buf(116));
  drc_bufs24211 : INVD5BWP7T port map(I => n_688, ZN => framebuffer_buf(41));
  drc_bufs24217 : INVD5BWP7T port map(I => n_694, ZN => framebuffer_buf(114));
  drc_bufs24223 : INVD5BWP7T port map(I => n_700, ZN => framebuffer_buf(113));
  drc_bufs24229 : INVD5BWP7T port map(I => n_706, ZN => framebuffer_buf(112));
  drc_bufs24235 : INVD5BWP7T port map(I => n_712, ZN => framebuffer_buf(107));
  drc_bufs24241 : INVD5BWP7T port map(I => n_718, ZN => framebuffer_buf(108));
  drc_bufs24247 : INVD5BWP7T port map(I => n_724, ZN => framebuffer_buf(42));
  drc_bufs24253 : INVD5BWP7T port map(I => n_730, ZN => framebuffer_buf(109));
  drc_bufs24259 : INVD5BWP7T port map(I => n_736, ZN => framebuffer_buf(110));
  drc_bufs24265 : INVD5BWP7T port map(I => n_742, ZN => framebuffer_buf(10));
  drc_bufs24271 : INVD5BWP7T port map(I => n_748, ZN => framebuffer_buf(43));
  drc_bufs24277 : INVD5BWP7T port map(I => n_754, ZN => framebuffer_buf(111));
  drc_bufs24283 : INVD5BWP7T port map(I => n_760, ZN => framebuffer_buf(44));
  drc_bufs24289 : INVD5BWP7T port map(I => n_766, ZN => framebuffer_buf(102));
  drc_bufs24295 : INVD5BWP7T port map(I => n_772, ZN => framebuffer_buf(101));
  drc_bufs24301 : INVD5BWP7T port map(I => n_778, ZN => framebuffer_buf(100));
  drc_bufs24307 : INVD5BWP7T port map(I => n_784, ZN => framebuffer_buf(99));
  drc_bufs24313 : INVD5BWP7T port map(I => n_790, ZN => framebuffer_buf(98));
  drc_bufs24319 : INVD5BWP7T port map(I => n_796, ZN => framebuffer_buf(97));
  drc_bufs24325 : INVD5BWP7T port map(I => n_802, ZN => framebuffer_buf(96));
  drc_bufs24331 : INVD5BWP7T port map(I => n_808, ZN => framebuffer_buf(45));
  drc_bufs24337 : INVD5BWP7T port map(I => n_814, ZN => framebuffer_buf(94));
  drc_bufs24343 : INVD5BWP7T port map(I => n_820, ZN => framebuffer_buf(93));
  drc_bufs24349 : INVD5BWP7T port map(I => n_826, ZN => framebuffer_buf(92));
  drc_bufs24355 : INVD5BWP7T port map(I => n_832, ZN => framebuffer_buf(115));
  drc_bufs24361 : INVD5BWP7T port map(I => n_838, ZN => framebuffer_buf(90));
  drc_bufs24367 : INVD5BWP7T port map(I => n_844, ZN => framebuffer_buf(89));
  drc_bufs24373 : INVD5BWP7T port map(I => n_850, ZN => framebuffer_buf(88));
  drc_bufs24379 : INVD5BWP7T port map(I => n_856, ZN => framebuffer_buf(46));
  drc_bufs24385 : INVD5BWP7T port map(I => n_862, ZN => framebuffer_buf(86));
  drc_bufs24391 : INVD5BWP7T port map(I => n_868, ZN => framebuffer_buf(85));
  drc_bufs24397 : INVD5BWP7T port map(I => n_874, ZN => framebuffer_buf(84));
  drc_bufs24403 : INVD5BWP7T port map(I => n_880, ZN => framebuffer_buf(11));
  drc_bufs24409 : INVD5BWP7T port map(I => n_886, ZN => framebuffer_buf(82));
  drc_bufs24415 : INVD5BWP7T port map(I => n_892, ZN => framebuffer_buf(12));
  drc_bufs24421 : INVD5BWP7T port map(I => n_898, ZN => framebuffer_buf(80));
  drc_bufs24427 : INVD5BWP7T port map(I => n_904, ZN => framebuffer_buf(47));
  drc_bufs24433 : INVD5BWP7T port map(I => n_910, ZN => framebuffer_buf(78));
  drc_bufs24439 : INVD5BWP7T port map(I => n_916, ZN => framebuffer_buf(77));
  drc_bufs24445 : INVD5BWP7T port map(I => n_922, ZN => framebuffer_buf(76));
  drc_bufs24451 : INVD5BWP7T port map(I => n_928, ZN => framebuffer_buf(119));
  drc_bufs24457 : INVD5BWP7T port map(I => n_934, ZN => framebuffer_buf(74));
  drc_bufs24463 : INVD5BWP7T port map(I => n_940, ZN => framebuffer_buf(48));
  drc_bufs24469 : INVD5BWP7T port map(I => n_946, ZN => framebuffer_buf(72));
  drc_bufs24475 : INVD5BWP7T port map(I => n_952, ZN => framebuffer_buf(49));
  drc_bufs24481 : INVD5BWP7T port map(I => n_958, ZN => framebuffer_buf(70));
  drc_bufs24487 : INVD5BWP7T port map(I => n_964, ZN => framebuffer_buf(69));
  drc_bufs24493 : INVD5BWP7T port map(I => n_970, ZN => framebuffer_buf(68));
  drc_bufs24499 : INVD5BWP7T port map(I => n_976, ZN => framebuffer_buf(123));
  drc_bufs24505 : INVD5BWP7T port map(I => n_982, ZN => framebuffer_buf(66));
  drc_bufs24511 : INVD5BWP7T port map(I => n_988, ZN => framebuffer_buf(155));
  drc_bufs24517 : INVD5BWP7T port map(I => n_994, ZN => framebuffer_buf(64));
  drc_bufs24523 : INVD5BWP7T port map(I => n_1000, ZN => framebuffer_buf(151));
  drc_bufs24529 : INVD5BWP7T port map(I => n_1006, ZN => framebuffer_buf(62));
  drc_bufs24535 : INVD5BWP7T port map(I => n_1012, ZN => framebuffer_buf(61));
  drc_bufs24541 : INVD5BWP7T port map(I => n_1018, ZN => framebuffer_buf(60));
  drc_bufs24547 : INVD5BWP7T port map(I => n_1024, ZN => framebuffer_buf(143));
  drc_bufs24553 : INVD5BWP7T port map(I => n_1030, ZN => framebuffer_buf(58));
  drc_bufs24559 : INVD5BWP7T port map(I => n_1036, ZN => framebuffer_buf(139));
  drc_bufs24565 : INVD5BWP7T port map(I => n_1042, ZN => framebuffer_buf(137));
  drc_bufs24571 : INVD5BWP7T port map(I => n_1048, ZN => framebuffer_buf(135));
  drc_bufs24577 : INVD5BWP7T port map(I => n_1054, ZN => framebuffer_buf(54));
  drc_bufs24583 : INVD5BWP7T port map(I => n_1060, ZN => framebuffer_buf(53));
  drc_bufs24589 : INVD5BWP7T port map(I => n_1066, ZN => framebuffer_buf(50));
  drc_bufs24595 : INVD5BWP7T port map(I => n_1072, ZN => framebuffer_buf(13));
  drc_bufs24601 : INVD5BWP7T port map(I => n_1078, ZN => framebuffer_buf(51));
  drc_bufs24607 : INVD5BWP7T port map(I => n_1084, ZN => framebuffer_buf(127));
  drc_bufs24613 : INVD5BWP7T port map(I => n_1090, ZN => framebuffer_buf(52));
  drc_bufs24619 : INVD5BWP7T port map(I => n_1096, ZN => framebuffer_buf(14));
  drc_bufs24625 : INVD5BWP7T port map(I => n_1102, ZN => framebuffer_buf(15));
  drc_bufs24631 : INVD5BWP7T port map(I => n_1108, ZN => framebuffer_buf(16));
  drc_bufs24637 : INVD5BWP7T port map(I => n_1114, ZN => framebuffer_buf(55));
  drc_bufs24643 : INVD5BWP7T port map(I => n_1120, ZN => framebuffer_buf(56));
  drc_bufs24649 : INVD5BWP7T port map(I => n_1126, ZN => framebuffer_buf(57));
  drc_bufs24655 : INVD5BWP7T port map(I => n_1132, ZN => framebuffer_buf(17));
  drc_bufs24661 : INVD5BWP7T port map(I => n_1138, ZN => framebuffer_buf(59));
  drc_bufs24667 : INVD5BWP7T port map(I => n_1144, ZN => framebuffer_buf(18));
  drc_bufs24673 : INVD5BWP7T port map(I => n_1150, ZN => framebuffer_buf(38));
  drc_bufs24679 : INVD5BWP7T port map(I => n_1156, ZN => framebuffer_buf(37));
  drc_bufs24685 : INVD5BWP7T port map(I => n_1162, ZN => framebuffer_buf(36));
  drc_bufs24691 : INVD5BWP7T port map(I => n_1168, ZN => framebuffer_buf(95));
  drc_bufs24697 : INVD5BWP7T port map(I => n_1174, ZN => framebuffer_buf(34));
  drc_bufs24703 : INVD5BWP7T port map(I => n_1180, ZN => framebuffer_buf(91));
  drc_bufs24709 : INVD5BWP7T port map(I => n_1186, ZN => framebuffer_buf(32));
  drc_bufs24715 : INVD5BWP7T port map(I => n_1192, ZN => framebuffer_buf(87));
  drc_bufs24721 : INVD5BWP7T port map(I => n_1198, ZN => framebuffer_buf(30));
  drc_bufs24727 : INVD5BWP7T port map(I => n_1204, ZN => framebuffer_buf(83));
  drc_bufs24733 : INVD5BWP7T port map(I => n_1210, ZN => framebuffer_buf(81));
  drc_bufs24739 : INVD5BWP7T port map(I => n_1216, ZN => framebuffer_buf(79));
  drc_bufs24745 : INVD5BWP7T port map(I => n_1222, ZN => framebuffer_buf(26));
  drc_bufs24751 : INVD5BWP7T port map(I => n_1228, ZN => framebuffer_buf(75));
  drc_bufs24757 : INVD5BWP7T port map(I => n_1234, ZN => framebuffer_buf(73));
  drc_bufs24763 : INVD5BWP7T port map(I => n_1240, ZN => framebuffer_buf(71));
  drc_bufs24769 : INVD5BWP7T port map(I => n_1246, ZN => framebuffer_buf(22));
  drc_bufs24775 : INVD5BWP7T port map(I => n_1252, ZN => framebuffer_buf(67));
  drc_bufs24781 : INVD5BWP7T port map(I => n_1258, ZN => framebuffer_buf(19));
  drc_bufs24787 : INVD5BWP7T port map(I => n_1264, ZN => framebuffer_buf(20));
  drc_bufs24793 : INVD5BWP7T port map(I => n_1270, ZN => framebuffer_buf(63));
  drc_bufs24799 : INVD5BWP7T port map(I => n_1276, ZN => framebuffer_buf(65));
  drc_bufs24805 : INVD5BWP7T port map(I => n_1282, ZN => framebuffer_buf(21));
  drc_bufs24811 : INVD5BWP7T port map(I => n_1288, ZN => framebuffer_buf(1));
  drc_bufs24817 : INVD5BWP7T port map(I => n_1294, ZN => framebuffer_buf(2));
  drc_bufs24823 : INVD5BWP7T port map(I => n_1300, ZN => framebuffer_buf(23));
  drc_bufs24829 : INVD5BWP7T port map(I => n_1306, ZN => framebuffer_buf(24));
  drc_bufs24835 : INVD5BWP7T port map(I => n_1312, ZN => framebuffer_buf(25));
  drc_bufs24841 : INVD5BWP7T port map(I => n_1318, ZN => framebuffer_buf(27));
  drc_bufs24847 : INVD5BWP7T port map(I => n_1324, ZN => framebuffer_buf(28));
  drc_bufs24853 : INVD5BWP7T port map(I => n_1330, ZN => framebuffer_buf(29));
  drc_bufs24859 : INVD5BWP7T port map(I => n_1336, ZN => framebuffer_buf(3));
  drc_bufs24865 : INVD5BWP7T port map(I => n_1342, ZN => framebuffer_buf(6));
  drc_bufs24871 : INVD5BWP7T port map(I => n_1348, ZN => framebuffer_buf(35));
  drc_bufs24877 : INVD5BWP7T port map(I => n_1354, ZN => framebuffer_buf(4));
  drc_bufs24883 : INVD5BWP7T port map(I => n_1362, ZN => framebuffer_buf(31));
  drc_bufs24889 : INVD5BWP7T port map(I => n_1368, ZN => framebuffer_buf(33));
  drc_bufs24895 : INVD5BWP7T port map(I => n_1374, ZN => framebuffer_buf(5));
  drc_bufs24901 : INVD5BWP7T port map(I => n_1380, ZN => calc_buf_out(23));
  drc_bufs24907 : INVD5BWP7T port map(I => n_1386, ZN => calc_buf_out(6));
  drc_bufs24913 : INVD5BWP7T port map(I => n_1392, ZN => calc_buf_out(9));
  drc_bufs24919 : INVD5BWP7T port map(I => n_1398, ZN => calc_buf_out(21));
  drc_bufs24925 : INVD5BWP7T port map(I => n_1404, ZN => calc_buf_out(1));
  drc_bufs24931 : INVD5BWP7T port map(I => n_1410, ZN => calc_buf_out(20));
  drc_bufs24937 : INVD5BWP7T port map(I => n_1416, ZN => calc_buf_out(12));
  drc_bufs24943 : INVD5BWP7T port map(I => n_1422, ZN => calc_buf_out(5));
  drc_bufs24949 : INVD5BWP7T port map(I => n_1428, ZN => calc_buf_out(15));
  drc_bufs24955 : INVD5BWP7T port map(I => n_1434, ZN => calc_buf_out(17));
  drc_bufs24961 : INVD5BWP7T port map(I => n_1440, ZN => calc_buf_out(16));
  drc_bufs24967 : INVD5BWP7T port map(I => n_1446, ZN => calc_buf_out(4));
  drc_bufs24973 : INVD5BWP7T port map(I => n_1452, ZN => calc_buf_out(10));
  drc_bufs24979 : INVD5BWP7T port map(I => n_1458, ZN => calc_buf_out(22));
  drc_bufs24985 : INVD5BWP7T port map(I => n_1464, ZN => calc_buf_out(8));
  drc_bufs24991 : INVD5BWP7T port map(I => n_1470, ZN => calc_buf_out(18));
  drc_bufs24997 : INVD5BWP7T port map(I => n_1476, ZN => calc_buf_out(0));
  drc_bufs25003 : INVD5BWP7T port map(I => n_1482, ZN => calc_buf_out(14));
  drc_bufs25009 : INVD5BWP7T port map(I => n_1488, ZN => calc_buf_out(2));
  drc_bufs25015 : INVD5BWP7T port map(I => n_1494, ZN => calc_buf_out(7));
  drc_bufs25021 : INVD5BWP7T port map(I => n_1500, ZN => calc_buf_out(19));
  drc_bufs25027 : INVD5BWP7T port map(I => n_1506, ZN => calc_buf_out(13));
  drc_bufs25033 : INVD5BWP7T port map(I => n_1512, ZN => calc_buf_out(11));
  drc_bufs25039 : INVD5BWP7T port map(I => n_1518, ZN => calc_buf_out(3));
  counter_reg_7 : DFKCND1BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => new_counter(7), Q => counter(7), QN => n_0);
  counter_reg_4 : DFKCND1BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => new_counter(4), Q => counter(4), QN => n_45);
  counter_reg_0 : DFKCND1BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => new_counter(0), Q => counter(0), QN => n_22);
  counter_reg_5 : DFKCND1BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => new_counter(5), Q => counter(5), QN => n_145);
  framebuffer_buf_reg_0 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_240, Q => framebuffer_buf_0_2288, QN => n_430);
  framebuffer_buf_reg_157 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_264, Q => framebuffer_buf_157_2445, QN => n_436);
  framebuffer_buf_reg_156 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_266, Q => framebuffer_buf_156_2444, QN => n_442);
  framebuffer_buf_reg_7 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_197, Q => framebuffer_buf_7_2295, QN => n_448);
  framebuffer_buf_reg_154 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_267, Q => framebuffer_buf_154_2442, QN => n_454);
  framebuffer_buf_reg_153 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_268, Q => framebuffer_buf_153_2441, QN => n_460);
  framebuffer_buf_reg_152 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_272, Q => framebuffer_buf_152_2440, QN => n_466);
  framebuffer_buf_reg_8 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_354, Q => framebuffer_buf_8_2296, QN => n_472);
  framebuffer_buf_reg_150 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_185, Q => FE_PHN184_framebuffer_buf_150_2438, QN => n_478);
  framebuffer_buf_reg_149 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_238, Q => framebuffer_buf_149_2437, QN => n_484);
  framebuffer_buf_reg_148 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_242, Q => framebuffer_buf_148_2436, QN => n_490);
  framebuffer_buf_reg_147 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_244, Q => framebuffer_buf_147_2435, QN => n_496);
  framebuffer_buf_reg_146 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_157, Q => framebuffer_buf_146_2434, QN => n_502);
  framebuffer_buf_reg_145 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_252, Q => framebuffer_buf_145_2433, QN => n_508);
  framebuffer_buf_reg_144 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_258, Q => framebuffer_buf_144_2432, QN => n_514);
  framebuffer_buf_reg_9 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_352, Q => framebuffer_buf_9_2297, QN => n_520);
  framebuffer_buf_reg_142 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_359, Q => FE_PHN87_framebuffer_buf_142_2430, QN => n_526);
  framebuffer_buf_reg_141 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_360, Q => framebuffer_buf_141_2429, QN => n_532);
  framebuffer_buf_reg_140 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_361, Q => framebuffer_buf_140_2428, QN => n_538);
  framebuffer_buf_reg_39 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_321, Q => framebuffer_buf_39_2327, QN => n_544);
  framebuffer_buf_reg_138 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_364, Q => FE_PHN155_framebuffer_buf_138_2426, QN => n_550);
  framebuffer_buf_reg_40 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_312, Q => framebuffer_buf_40_2328, QN => n_556);
  framebuffer_buf_reg_136 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_371, Q => FE_PHN161_framebuffer_buf_136_2424, QN => n_562);
  framebuffer_buf_reg_103 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_178, Q => framebuffer_buf_103_2391, QN => n_568);
  framebuffer_buf_reg_134 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_194, Q => framebuffer_buf_134_2422, QN => n_574);
  framebuffer_buf_reg_133 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_256, Q => framebuffer_buf_133_2421, QN => n_580);
  framebuffer_buf_reg_132 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_265, Q => framebuffer_buf_132_2420, QN => n_586);
  framebuffer_buf_reg_131 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_269, Q => framebuffer_buf_131_2419, QN => n_592);
  framebuffer_buf_reg_130 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_273, Q => FE_PHN167_framebuffer_buf_130_2418, QN => n_598);
  framebuffer_buf_reg_129 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_274, Q => framebuffer_buf_129_2417, QN => n_604);
  framebuffer_buf_reg_128 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_277, Q => FE_PHN51_framebuffer_buf_128_2416, QN => n_610);
  framebuffer_buf_reg_104 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_172, Q => FE_PHN187_framebuffer_buf_104_2392, QN => n_616);
  framebuffer_buf_reg_126 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_340, Q => framebuffer_buf_126_2414, QN => n_622);
  framebuffer_buf_reg_125 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_249, Q => framebuffer_buf_125_2413, QN => n_628);
  framebuffer_buf_reg_124 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_158, Q => framebuffer_buf_124_2412, QN => n_634);
  framebuffer_buf_reg_105 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_171, Q => framebuffer_buf_105_2393, QN => n_640);
  framebuffer_buf_reg_122 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_160, Q => framebuffer_buf_122_2410, QN => n_646);
  framebuffer_buf_reg_121 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_161, Q => framebuffer_buf_121_2409, QN => n_652);
  framebuffer_buf_reg_120 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_162, Q => framebuffer_buf_120_2408, QN => n_658);
  framebuffer_buf_reg_106 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_168, Q => framebuffer_buf_106_2394, QN => n_664);
  framebuffer_buf_reg_118 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_292, Q => framebuffer_buf_118_2406, QN => n_670);
  framebuffer_buf_reg_117 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_293, Q => framebuffer_buf_117_2405, QN => n_676);
  framebuffer_buf_reg_116 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_297, Q => framebuffer_buf_116_2404, QN => n_682);
  framebuffer_buf_reg_41 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_234, Q => framebuffer_buf_41_2329, QN => n_688);
  framebuffer_buf_reg_114 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_299, Q => framebuffer_buf_114_2402, QN => n_694);
  framebuffer_buf_reg_113 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_305, Q => framebuffer_buf_113_2401, QN => n_700);
  framebuffer_buf_reg_112 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_309, Q => framebuffer_buf_112_2400, QN => n_706);
  framebuffer_buf_reg_107 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_167, Q => framebuffer_buf_107_2395, QN => n_712);
  framebuffer_buf_reg_108 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_166, Q => framebuffer_buf_108_2396, QN => n_718);
  framebuffer_buf_reg_42 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_228, Q => framebuffer_buf_42_2330, QN => n_724);
  framebuffer_buf_reg_109 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_165, Q => FE_PHN175_framebuffer_buf_109_2397, QN => n_730);
  framebuffer_buf_reg_110 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => n_163, Q => framebuffer_buf_110_2398, QN => n_736);
  framebuffer_buf_reg_10 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_348, Q => framebuffer_buf_10_2298, QN => n_742);
  framebuffer_buf_reg_43 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_191, Q => framebuffer_buf_43_2331, QN => n_748);
  framebuffer_buf_reg_111 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_164, Q => framebuffer_buf_111_2399, QN => n_754);
  framebuffer_buf_reg_44 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_221, Q => FE_PHN171_framebuffer_buf_44_2332, QN => n_760);
  framebuffer_buf_reg_102 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_179, Q => framebuffer_buf_102_2390, QN => n_766);
  framebuffer_buf_reg_101 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_180, Q => framebuffer_buf_101_2389, QN => n_772);
  framebuffer_buf_reg_100 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_182, Q => framebuffer_buf_100_2388, QN => n_778);
  framebuffer_buf_reg_99 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_183, Q => FE_PHN134_framebuffer_buf_99_2387, QN => n_784);
  framebuffer_buf_reg_98 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_184, Q => FE_PHN98_framebuffer_buf_98_2386, QN => n_790);
  framebuffer_buf_reg_97 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_188, Q => framebuffer_buf_97_2385, QN => n_796);
  framebuffer_buf_reg_96 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_190, Q => framebuffer_buf_96_2384, QN => n_802);
  framebuffer_buf_reg_45 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_220, Q => framebuffer_buf_45_2333, QN => n_808);
  framebuffer_buf_reg_94 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_193, Q => framebuffer_buf_94_2382, QN => n_814);
  framebuffer_buf_reg_93 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => n_195, Q => framebuffer_buf_93_2381, QN => n_820);
  framebuffer_buf_reg_92 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_196, Q => framebuffer_buf_92_2380, QN => n_826);
  framebuffer_buf_reg_115 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_298, Q => framebuffer_buf_115_2403, QN => n_832);
  framebuffer_buf_reg_90 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => n_200, Q => framebuffer_buf_90_2378, QN => n_838);
  framebuffer_buf_reg_89 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => n_207, Q => framebuffer_buf_89_2377, QN => n_844);
  framebuffer_buf_reg_88 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => n_209, Q => framebuffer_buf_88_2376, QN => n_850);
  framebuffer_buf_reg_46 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_176, Q => framebuffer_buf_46_2334, QN => n_856);
  framebuffer_buf_reg_86 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_211, Q => framebuffer_buf_86_2374, QN => n_862);
  framebuffer_buf_reg_85 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_215, Q => framebuffer_buf_85_2373, QN => n_868);
  framebuffer_buf_reg_84 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_217, Q => framebuffer_buf_84_2372, QN => n_874);
  framebuffer_buf_reg_11 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_346, Q => framebuffer_buf_11_2299, QN => n_880);
  framebuffer_buf_reg_82 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_223, Q => FE_PHN5_framebuffer_buf_82_2370, QN => n_886);
  framebuffer_buf_reg_12 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_344, Q => FE_PHN122_framebuffer_buf_12_2300, QN => n_892);
  framebuffer_buf_reg_80 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_308, Q => framebuffer_buf_80_2368, QN => n_898);
  framebuffer_buf_reg_47 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_175, Q => FE_PHN135_framebuffer_buf_47_2335, QN => n_904);
  framebuffer_buf_reg_78 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_307, Q => FE_PHN148_framebuffer_buf_78_2366, QN => n_910);
  framebuffer_buf_reg_77 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => n_236, Q => framebuffer_buf_77_2365, QN => n_916);
  framebuffer_buf_reg_76 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => n_237, Q => framebuffer_buf_76_2364, QN => n_922);
  framebuffer_buf_reg_119 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_291, Q => framebuffer_buf_119_2407, QN => n_928);
  framebuffer_buf_reg_74 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => n_241, Q => framebuffer_buf_74_2362, QN => n_934);
  framebuffer_buf_reg_48 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_320, Q => framebuffer_buf_48_2336, QN => n_940);
  framebuffer_buf_reg_72 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => n_247, Q => framebuffer_buf_72_2360, QN => n_946);
  framebuffer_buf_reg_49 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_319, Q => framebuffer_buf_49_2337, QN => n_952);
  framebuffer_buf_reg_70 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => n_254, Q => framebuffer_buf_70_2358, QN => n_958);
  framebuffer_buf_reg_69 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => n_253, Q => framebuffer_buf_69_2357, QN => n_964);
  framebuffer_buf_reg_68 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => n_314, Q => framebuffer_buf_68_2356, QN => n_970);
  framebuffer_buf_reg_123 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_159, Q => framebuffer_buf_123_2411, QN => n_976);
  framebuffer_buf_reg_66 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => n_259, Q => framebuffer_buf_66_2354, QN => n_982);
  framebuffer_buf_reg_155 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_295, Q => framebuffer_buf_155_2443, QN => n_988);
  framebuffer_buf_reg_64 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => n_263, Q => framebuffer_buf_64_2352, QN => n_994);
  framebuffer_buf_reg_151 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_181, Q => FE_PHN162_framebuffer_buf_151_2439, QN => n_1000);
  framebuffer_buf_reg_62 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_174, Q => framebuffer_buf_62_2350, QN => n_1006);
  framebuffer_buf_reg_61 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_198, Q => framebuffer_buf_61_2349, QN => n_1012);
  framebuffer_buf_reg_60 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_201, Q => framebuffer_buf_60_2348, QN => n_1018);
  framebuffer_buf_reg_143 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_358, Q => framebuffer_buf_143_2431, QN => n_1024);
  framebuffer_buf_reg_58 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_208, Q => framebuffer_buf_58_2346, QN => n_1030);
  framebuffer_buf_reg_139 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_363, Q => FE_PHN88_framebuffer_buf_139_2427, QN => n_1036);
  framebuffer_buf_reg_137 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_368, Q => FE_PHN99_framebuffer_buf_137_2425, QN => n_1042);
  framebuffer_buf_reg_135 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_323, Q => FE_PHN107_framebuffer_buf_135_2423, QN => n_1048);
  framebuffer_buf_reg_54 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_313, Q => framebuffer_buf_54_2342, QN => n_1054);
  framebuffer_buf_reg_53 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_255, Q => framebuffer_buf_53_2341, QN => n_1060);
  framebuffer_buf_reg_50 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_189, Q => framebuffer_buf_50_2338, QN => n_1066);
  framebuffer_buf_reg_13 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_342, Q => framebuffer_buf_13_2301, QN => n_1072);
  framebuffer_buf_reg_51 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_315, Q => framebuffer_buf_51_2339, QN => n_1078);
  framebuffer_buf_reg_127 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_338, Q => framebuffer_buf_127_2415, QN => n_1084);
  framebuffer_buf_reg_52 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_316, Q => framebuffer_buf_52_2340, QN => n_1090);
  framebuffer_buf_reg_14 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_334, Q => FE_PHN186_framebuffer_buf_14_2302, QN => n_1096);
  framebuffer_buf_reg_15 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_333, Q => framebuffer_buf_15_2303, QN => n_1102);
  framebuffer_buf_reg_16 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_177, Q => framebuffer_buf_16_2304, QN => n_1108);
  framebuffer_buf_reg_55 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_310, Q => framebuffer_buf_55_2343, QN => n_1114);
  framebuffer_buf_reg_56 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_218, Q => framebuffer_buf_56_2344, QN => n_1120);
  framebuffer_buf_reg_57 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_214, Q => framebuffer_buf_57_2345, QN => n_1126);
  framebuffer_buf_reg_17 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_306, Q => framebuffer_buf_17_2305, QN => n_1132);
  framebuffer_buf_reg_59 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_204, Q => FE_PHN106_framebuffer_buf_59_2347, QN => n_1138);
  framebuffer_buf_reg_18 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_302, Q => framebuffer_buf_18_2306, QN => n_1144);
  framebuffer_buf_reg_38 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_322, Q => framebuffer_buf_38_2326, QN => n_1150);
  framebuffer_buf_reg_37 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_332, Q => framebuffer_buf_37_2325, QN => n_1156);
  framebuffer_buf_reg_36 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_325, Q => framebuffer_buf_36_2324, QN => n_1162);
  framebuffer_buf_reg_95 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_192, Q => framebuffer_buf_95_2383, QN => n_1168);
  framebuffer_buf_reg_34 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_326, Q => framebuffer_buf_34_2322, QN => n_1174);
  framebuffer_buf_reg_91 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_199, Q => framebuffer_buf_91_2379, QN => n_1180);
  framebuffer_buf_reg_32 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_331, Q => FE_PHN147_framebuffer_buf_32_2320, QN => n_1186);
  framebuffer_buf_reg_87 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_210, Q => framebuffer_buf_87_2375, QN => n_1192);
  framebuffer_buf_reg_30 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_279, Q => framebuffer_buf_30_2318, QN => n_1198);
  framebuffer_buf_reg_83 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_219, Q => framebuffer_buf_83_2371, QN => n_1204);
  framebuffer_buf_reg_81 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_226, Q => framebuffer_buf_81_2369, QN => n_1210);
  framebuffer_buf_reg_79 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_235, Q => framebuffer_buf_79_2367, QN => n_1216);
  framebuffer_buf_reg_26 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_283, Q => framebuffer_buf_26_2314, QN => n_1222);
  framebuffer_buf_reg_75 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_239, Q => framebuffer_buf_75_2363, QN => n_1228);
  framebuffer_buf_reg_73 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_243, Q => framebuffer_buf_73_2361, QN => n_1234);
  framebuffer_buf_reg_71 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => n_248, Q => framebuffer_buf_71_2359, QN => n_1240);
  framebuffer_buf_reg_22 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_289, Q => framebuffer_buf_22_2310, QN => n_1246);
  framebuffer_buf_reg_67 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_257, Q => framebuffer_buf_67_2355, QN => n_1252);
  framebuffer_buf_reg_19 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_296, Q => framebuffer_buf_19_2307, QN => n_1258);
  framebuffer_buf_reg_20 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_294, Q => framebuffer_buf_20_2308, QN => n_1264);
  framebuffer_buf_reg_63 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_173, Q => framebuffer_buf_63_2351, QN => n_1270);
  framebuffer_buf_reg_65 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_13, D => n_260, Q => framebuffer_buf_65_2353, QN => n_1276);
  framebuffer_buf_reg_21 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_290, Q => framebuffer_buf_21_2309, QN => n_1282);
  framebuffer_buf_reg_1 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_231, Q => framebuffer_buf_1_2289, QN => n_1288);
  framebuffer_buf_reg_2 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_227, Q => framebuffer_buf_2_2290, QN => n_1294);
  framebuffer_buf_reg_23 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_288, Q => framebuffer_buf_23_2311, QN => n_1300);
  framebuffer_buf_reg_24 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_287, Q => framebuffer_buf_24_2312, QN => n_1306);
  framebuffer_buf_reg_25 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_286, Q => framebuffer_buf_25_2313, QN => n_1312);
  framebuffer_buf_reg_27 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_282, Q => framebuffer_buf_27_2315, QN => n_1318);
  framebuffer_buf_reg_28 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_281, Q => framebuffer_buf_28_2316, QN => n_1324);
  framebuffer_buf_reg_29 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_280, Q => framebuffer_buf_29_2317, QN => n_1330);
  framebuffer_buf_reg_3 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_222, Q => FE_PHN121_framebuffer_buf_3_2291, QN => n_1336);
  framebuffer_buf_reg_6 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_202, Q => framebuffer_buf_6_2294, QN => n_1342);
  framebuffer_buf_reg_35 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_324, Q => framebuffer_buf_35_2323, QN => n_1348);
  framebuffer_buf_reg_4 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_216, Q => FE_PHN50_framebuffer_buf_4_2292, QN => n_1354);
  framebuffer_buf_reg_31 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_278, Q => framebuffer_buf_31_2319, QN => n_1362);
  framebuffer_buf_reg_33 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_328, Q => framebuffer_buf_33_2321, QN => n_1368);
  framebuffer_buf_reg_5 : DFKCND0BWP7T port map(CN => FE_OFN1_FE_DBTN0_reset, CP => CTS_13, D => n_203, Q => framebuffer_buf_5_2293, QN => n_1374);
  calc_buf_out_reg_23 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_365, Q => calc_buf_out_23_2287, QN => n_1380);
  calc_buf_out_reg_6 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => new_calc_buf_out(6), Q => calc_buf_out_6_2270, QN => n_1386);
  calc_buf_out_reg_9 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_386, Q => calc_buf_out_9_2273, QN => n_1392);
  calc_buf_out_reg_21 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_370, Q => calc_buf_out_21_2285, QN => n_1398);
  calc_buf_out_reg_1 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => new_calc_buf_out(1), Q => calc_buf_out_1_2265, QN => n_1404);
  calc_buf_out_reg_20 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_355, Q => calc_buf_out_20_2284, QN => n_1410);
  calc_buf_out_reg_12 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_381, Q => FE_PHN93_calc_buf_out_12_2276, QN => n_1416);
  calc_buf_out_reg_5 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => new_calc_buf_out(5), Q => calc_buf_out_5_2269, QN => n_1422);
  calc_buf_out_reg_15 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_379, Q => calc_buf_out_15_2279, QN => n_1428);
  calc_buf_out_reg_17 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_375, Q => FE_PHN23_calc_buf_out_17_2281, QN => n_1434);
  calc_buf_out_reg_16 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_378, Q => FE_PHN41_calc_buf_out_16_2280, QN => n_1440);
  calc_buf_out_reg_4 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => new_calc_buf_out(4), Q => calc_buf_out_4_2268, QN => n_1446);
  calc_buf_out_reg_10 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_383, Q => calc_buf_out_10_2274, QN => n_1452);
  calc_buf_out_reg_22 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_369, Q => FE_PHN28_calc_buf_out_22_2286, QN => n_1458);
  calc_buf_out_reg_8 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_387, Q => calc_buf_out_8_2272, QN => n_1464);
  calc_buf_out_reg_18 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_374, Q => calc_buf_out_18_2282, QN => n_1470);
  calc_buf_out_reg_0 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => new_calc_buf_out(0), Q => calc_buf_out_0_2264, QN => n_1476);
  calc_buf_out_reg_14 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_380, Q => calc_buf_out_14_2278, QN => n_1482);
  calc_buf_out_reg_2 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => new_calc_buf_out(2), Q => calc_buf_out_2_2266, QN => n_1488);
  calc_buf_out_reg_7 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => new_calc_buf_out(7), Q => calc_buf_out_7_2271, QN => n_1494);
  calc_buf_out_reg_19 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => n_394, Q => calc_buf_out_19_2283, QN => n_1500);
  calc_buf_out_reg_13 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_362, Q => FE_PHN37_calc_buf_out_13_2277, QN => n_1506);
  calc_buf_out_reg_11 : DFKCND0BWP7T port map(CN => FE_OFN0_FE_DBTN0_reset, CP => CTS_12, D => n_382, Q => calc_buf_out_11_2275, QN => n_1512);
  calc_buf_out_reg_3 : DFKCND0BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_12, D => new_calc_buf_out(3), Q => calc_buf_out_3_2267, QN => n_1518);
  g2 : IND2D1BWP7T port map(A1 => n_83, B1 => counter(0), ZN => n_1522);
  g25416 : IND2D1BWP7T port map(A1 => n_69, B1 => n_76, ZN => n_1523);

end routed;
