library IEEE;
use IEEE.std_logic_1164.ALL;

entity sqi_controller_tb is
end sqi_controller_tb;

