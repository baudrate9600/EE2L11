configuration sram_interface_routed_cfg of sram_interface is
   for routed
   end for;
end sram_interface_routed_cfg;
