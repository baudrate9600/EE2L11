library IEEE;
use IEEE.std_logic_1164.ALL;

entity sram_interface_tb is
end sram_interface_tb;

