configuration sqi_synthesised_cfg of sqi is
   for synthesised
   end for;
end sqi_synthesised_cfg;
