library IEEE;
use IEEE.std_logic_1164.ALL;

entity sqi_tb is
end sqi_tb;

