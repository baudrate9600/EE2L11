configuration gen25mhz_behaviour_cfg of gen25mhz is
   for behaviour
   end for;
end gen25mhz_behaviour_cfg;
