configuration prescaler_behaviour_cfg of prescaler is
   for behaviour
   end for;
end prescaler_behaviour_cfg;
