library IEEE;
use IEEE.std_logic_1164.ALL;

entity line_buffer_tb is
end line_buffer_tb;

