
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture synthesised of memory is

  component DFKCNQD1BWP7T
    port(CP, CN, D : in std_logic; Q : out std_logic);
  end component;

  component LHQD1BWP7T
    port(E, D : in std_logic; Q : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component IOA21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component IIND4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component CKND4BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component LHD1BWP7T
    port(E, D : in std_logic; Q, QN : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component DFXQD1BWP7T
    port(CP, DA, DB, SA : in std_logic; Q : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IND3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component CKAN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component CKND0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component ND2D4BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INVD4BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CP, CN, D : in std_logic; Q, QN : out std_logic);
  end component;

  component EDFD0BWP7T
    port(CP, D, E : in std_logic; Q, QN : out std_logic);
  end component;

  signal new_counter : std_logic_vector(7 downto 0);
  signal counter : std_logic_vector(7 downto 0);
  signal new_calc_buf_out : std_logic_vector(23 downto 0);
  signal state : std_logic_vector(3 downto 0);
  signal new_framebuffer_buf : std_logic_vector(157 downto 0);
  signal new_row_buf : std_logic_vector(5 downto 0);
  signal row_buf : std_logic_vector(5 downto 0);
  signal UNCONNECTED, UNCONNECTED0, UNCONNECTED1, UNCONNECTED2, UNCONNECTED3 : std_logic;
  signal UNCONNECTED4, UNCONNECTED5, UNCONNECTED6, calc_buf_out_0_3514, calc_buf_out_1_3515 : std_logic;
  signal calc_buf_out_2_3516, calc_buf_out_3_3517, calc_buf_out_4_3518, calc_buf_out_5_3519, calc_buf_out_6_3520 : std_logic;
  signal calc_buf_out_7_3521, calc_buf_out_8_3522, calc_buf_out_9_3523, calc_buf_out_10_3524, calc_buf_out_11_3525 : std_logic;
  signal calc_buf_out_12_3526, calc_buf_out_13_3527, calc_buf_out_14_3528, calc_buf_out_15_3529, calc_buf_out_16_3530 : std_logic;
  signal calc_buf_out_17_3531, calc_buf_out_18_3532, calc_buf_out_19_3533, calc_buf_out_20_3534, calc_buf_out_21_3535 : std_logic;
  signal calc_buf_out_22_3536, calc_buf_out_23_3537, framebuffer_buf_0_3538, framebuffer_buf_1_3539, framebuffer_buf_2_3540 : std_logic;
  signal framebuffer_buf_3_3541, framebuffer_buf_4_3542, framebuffer_buf_5_3543, framebuffer_buf_6_3544, framebuffer_buf_7_3545 : std_logic;
  signal framebuffer_buf_8_3546, framebuffer_buf_9_3547, framebuffer_buf_10_3548, framebuffer_buf_11_3549, framebuffer_buf_12_3550 : std_logic;
  signal framebuffer_buf_13_3551, framebuffer_buf_14_3552, framebuffer_buf_15_3553, framebuffer_buf_16_3554, framebuffer_buf_17_3555 : std_logic;
  signal framebuffer_buf_18_3556, framebuffer_buf_19_3557, framebuffer_buf_20_3558, framebuffer_buf_21_3559, framebuffer_buf_22_3560 : std_logic;
  signal framebuffer_buf_23_3561, framebuffer_buf_24_3562, framebuffer_buf_25_3563, framebuffer_buf_26_3564, framebuffer_buf_27_3565 : std_logic;
  signal framebuffer_buf_28_3566, framebuffer_buf_29_3567, framebuffer_buf_30_3568, framebuffer_buf_31_3569, framebuffer_buf_32_3570 : std_logic;
  signal framebuffer_buf_33_3571, framebuffer_buf_34_3572, framebuffer_buf_35_3573, framebuffer_buf_36_3574, framebuffer_buf_37_3575 : std_logic;
  signal framebuffer_buf_38_3576, framebuffer_buf_39_3577, framebuffer_buf_40_3578, framebuffer_buf_41_3579, framebuffer_buf_42_3580 : std_logic;
  signal framebuffer_buf_43_3581, framebuffer_buf_44_3582, framebuffer_buf_45_3583, framebuffer_buf_46_3584, framebuffer_buf_47_3585 : std_logic;
  signal framebuffer_buf_48_3586, framebuffer_buf_49_3587, framebuffer_buf_50_3588, framebuffer_buf_51_3589, framebuffer_buf_52_3590 : std_logic;
  signal framebuffer_buf_53_3591, framebuffer_buf_54_3592, framebuffer_buf_55_3593, framebuffer_buf_56_3594, framebuffer_buf_57_3595 : std_logic;
  signal framebuffer_buf_58_3596, framebuffer_buf_59_3597, framebuffer_buf_60_3598, framebuffer_buf_61_3599, framebuffer_buf_62_3600 : std_logic;
  signal framebuffer_buf_63_3601, framebuffer_buf_64_3602, framebuffer_buf_65_3603, framebuffer_buf_66_3604, framebuffer_buf_67_3605 : std_logic;
  signal framebuffer_buf_68_3606, framebuffer_buf_69_3607, framebuffer_buf_70_3608, framebuffer_buf_71_3609, framebuffer_buf_72_3610 : std_logic;
  signal framebuffer_buf_73_3611, framebuffer_buf_74_3612, framebuffer_buf_75_3613, framebuffer_buf_76_3614, framebuffer_buf_77_3615 : std_logic;
  signal framebuffer_buf_78_3616, framebuffer_buf_79_3617, framebuffer_buf_80_3618, framebuffer_buf_81_3619, framebuffer_buf_82_3620 : std_logic;
  signal framebuffer_buf_83_3621, framebuffer_buf_84_3622, framebuffer_buf_85_3623, framebuffer_buf_86_3624, framebuffer_buf_87_3625 : std_logic;
  signal framebuffer_buf_88_3626, framebuffer_buf_89_3627, framebuffer_buf_90_3628, framebuffer_buf_91_3629, framebuffer_buf_92_3630 : std_logic;
  signal framebuffer_buf_93_3631, framebuffer_buf_94_3632, framebuffer_buf_95_3633, framebuffer_buf_96_3634, framebuffer_buf_97_3635 : std_logic;
  signal framebuffer_buf_98_3636, framebuffer_buf_99_3637, framebuffer_buf_100_3638, framebuffer_buf_101_3639, framebuffer_buf_102_3640 : std_logic;
  signal framebuffer_buf_103_3641, framebuffer_buf_104_3642, framebuffer_buf_105_3643, framebuffer_buf_106_3644, framebuffer_buf_107_3645 : std_logic;
  signal framebuffer_buf_108_3646, framebuffer_buf_109_3647, framebuffer_buf_110_3648, framebuffer_buf_111_3649, framebuffer_buf_112_3650 : std_logic;
  signal framebuffer_buf_113_3651, framebuffer_buf_114_3652, framebuffer_buf_115_3653, framebuffer_buf_116_3654, framebuffer_buf_117_3655 : std_logic;
  signal framebuffer_buf_118_3656, framebuffer_buf_119_3657, framebuffer_buf_120_3658, framebuffer_buf_121_3659, framebuffer_buf_122_3660 : std_logic;
  signal framebuffer_buf_123_3661, framebuffer_buf_124_3662, framebuffer_buf_125_3663, framebuffer_buf_126_3664, framebuffer_buf_127_3665 : std_logic;
  signal framebuffer_buf_128_3666, framebuffer_buf_129_3667, framebuffer_buf_130_3668, framebuffer_buf_131_3669, framebuffer_buf_132_3670 : std_logic;
  signal framebuffer_buf_133_3671, framebuffer_buf_134_3672, framebuffer_buf_135_3673, framebuffer_buf_136_3674, framebuffer_buf_137_3675 : std_logic;
  signal framebuffer_buf_138_3676, framebuffer_buf_139_3677, framebuffer_buf_140_3678, framebuffer_buf_141_3679, framebuffer_buf_142_3680 : std_logic;
  signal framebuffer_buf_143_3681, framebuffer_buf_144_3682, framebuffer_buf_145_3683, framebuffer_buf_146_3684, framebuffer_buf_147_3685 : std_logic;
  signal framebuffer_buf_148_3686, framebuffer_buf_149_3687, framebuffer_buf_150_3688, framebuffer_buf_151_3689, framebuffer_buf_152_3690 : std_logic;
  signal framebuffer_buf_153_3691, framebuffer_buf_154_3692, framebuffer_buf_155_3693, framebuffer_buf_156_3694, framebuffer_buf_157_3695 : std_logic;
  signal n_1, n_2, n_3, n_4, n_5 : std_logic;
  signal n_6, n_7, n_8, n_9, n_10 : std_logic;
  signal n_11, n_12, n_13, n_14, n_16 : std_logic;
  signal n_17, n_18, n_19, n_20, n_21 : std_logic;
  signal n_22, n_23, n_24, n_25, n_26 : std_logic;
  signal n_28, n_29, n_30, n_32, n_33 : std_logic;
  signal n_34, n_35, n_36, n_37, n_38 : std_logic;
  signal n_39, n_40, n_41, n_42, n_43 : std_logic;
  signal n_44, n_45, n_46, n_47, n_48 : std_logic;
  signal n_49, n_50, n_51, n_52, n_53 : std_logic;
  signal n_54, n_55, n_56, n_57, n_59 : std_logic;
  signal n_60, n_61, n_62, n_63, n_64 : std_logic;
  signal n_65, n_66, n_67, n_68, n_69 : std_logic;
  signal n_70, n_71, n_72, n_73, n_74 : std_logic;
  signal n_75, n_76, n_77, n_78, n_79 : std_logic;
  signal n_80, n_81, n_82, n_83, n_84 : std_logic;
  signal n_85, n_86, n_87, n_88, n_89 : std_logic;
  signal n_90, n_91, n_92, n_93, n_94 : std_logic;
  signal n_95, n_96, n_97, n_98, n_99 : std_logic;
  signal n_100, n_101, n_102, n_103, n_104 : std_logic;
  signal n_105, n_106, n_107, n_108, n_109 : std_logic;
  signal n_110, n_111, n_112, n_113, n_114 : std_logic;
  signal n_115, n_116, n_117, n_118, n_119 : std_logic;
  signal n_120, n_122, n_123, n_124, n_125 : std_logic;
  signal n_126, n_127, n_128, n_129, n_130 : std_logic;
  signal n_131, n_132, n_133, n_134, n_135 : std_logic;
  signal n_136, n_137, n_138, n_139, n_140 : std_logic;
  signal n_141, n_142, n_143, n_144, n_145 : std_logic;
  signal n_146, n_147, n_148, n_149, n_150 : std_logic;
  signal n_151, n_152, n_153, n_154, n_155 : std_logic;
  signal n_156, n_157, n_158, n_159, n_160 : std_logic;
  signal n_161, n_162, n_163, n_164, n_165 : std_logic;
  signal n_166, n_167, n_168, n_169, n_170 : std_logic;
  signal n_171, n_172, n_173, n_174, n_175 : std_logic;
  signal n_176, n_177, n_178, n_179, n_180 : std_logic;
  signal n_181, n_182, n_183, n_184, n_185 : std_logic;
  signal n_186, n_187, n_188, n_189, n_190 : std_logic;
  signal n_191, n_192, n_193, n_194, n_195 : std_logic;
  signal n_196, n_197, n_198, n_199, n_200 : std_logic;
  signal n_201, n_202, n_203, n_204, n_205 : std_logic;
  signal n_206, n_207, n_208, n_209, n_210 : std_logic;
  signal n_211, n_212, n_213, n_214, n_215 : std_logic;
  signal n_216, n_217, n_218, n_219, n_220 : std_logic;
  signal n_221, n_222, n_223, n_224, n_225 : std_logic;
  signal n_226, n_227, n_228, n_229, n_230 : std_logic;
  signal n_231, n_239, n_240, n_241, n_242 : std_logic;
  signal n_243, n_244, n_245, n_246, n_247 : std_logic;
  signal n_248, n_249, n_250, n_251, n_252 : std_logic;
  signal n_253, n_254, n_255, n_256, n_257 : std_logic;
  signal n_258, n_259, n_260, n_261, n_262 : std_logic;
  signal n_263, n_264, n_265, n_266, n_267 : std_logic;
  signal n_268, n_269, n_270, n_271, n_272 : std_logic;
  signal n_273, n_274, n_276, n_277, n_278 : std_logic;
  signal n_279, n_280, n_281, n_282, n_283 : std_logic;
  signal n_284, n_285, n_286, n_287, n_288 : std_logic;
  signal n_289, n_290, n_291, n_292, n_293 : std_logic;
  signal n_294, n_296, n_297, n_298, n_299 : std_logic;
  signal n_300, n_301, n_302, n_304, n_305 : std_logic;
  signal n_306, n_307, n_308, n_309, n_310 : std_logic;
  signal n_311, n_312, n_313, n_314, n_315 : std_logic;
  signal n_316, n_317, n_318, n_319, n_321 : std_logic;
  signal n_322, n_323, n_324, n_325, n_326 : std_logic;
  signal n_327, n_328, n_329, n_330, n_331 : std_logic;
  signal n_332, n_333, n_334, n_335, n_336 : std_logic;
  signal n_337, n_338, n_339, n_340, n_341 : std_logic;
  signal n_342, n_343, n_344, n_345, n_346 : std_logic;
  signal n_347, n_349, n_350, n_351, n_352 : std_logic;
  signal n_353, n_354, n_355, n_356, n_357 : std_logic;
  signal n_360, n_362, n_363, n_364, n_365 : std_logic;
  signal n_366, n_367, n_368, n_369, n_389 : std_logic;
  signal n_392, n_398, n_404, n_410, n_416 : std_logic;
  signal n_422, n_428, n_434, n_440, n_446 : std_logic;
  signal n_452, n_458, n_464, n_470, n_476 : std_logic;
  signal n_482, n_488, n_494, n_500, n_506 : std_logic;
  signal n_512, n_518, n_524, n_530, n_536 : std_logic;
  signal n_542, n_548, n_554, n_560, n_566 : std_logic;
  signal n_572, n_578, n_584, n_590, n_596 : std_logic;
  signal n_602, n_608, n_614, n_620, n_626 : std_logic;
  signal n_632, n_638, n_644, n_650, n_656 : std_logic;
  signal n_662, n_668, n_674, n_680, n_686 : std_logic;
  signal n_692, n_698, n_704, n_710, n_716 : std_logic;
  signal n_722, n_728, n_734, n_740, n_746 : std_logic;
  signal n_752, n_758, n_764, n_770, n_776 : std_logic;
  signal n_782, n_788, n_794, n_800, n_806 : std_logic;
  signal n_812, n_818, n_824, n_830, n_836 : std_logic;
  signal n_842, n_848, n_854, n_860, n_866 : std_logic;
  signal n_872, n_878, n_884, n_890, n_896 : std_logic;
  signal n_902, n_908, n_914, n_920, n_926 : std_logic;
  signal n_932, n_938, n_944, n_950, n_956 : std_logic;
  signal n_962, n_968, n_974, n_980, n_986 : std_logic;
  signal n_992, n_998, n_1004, n_1010, n_1016 : std_logic;
  signal n_1022, n_1028, n_1034, n_1040, n_1046 : std_logic;
  signal n_1052, n_1058, n_1064, n_1070, n_1076 : std_logic;
  signal n_1082, n_1088, n_1094, n_1100, n_1106 : std_logic;
  signal n_1112, n_1118, n_1124, n_1130, n_1136 : std_logic;
  signal n_1142, n_1148, n_1154, n_1160, n_1166 : std_logic;
  signal n_1172, n_1178, n_1184, n_1190, n_1196 : std_logic;
  signal n_1202, n_1208, n_1214, n_1220, n_1226 : std_logic;
  signal n_1232, n_1238, n_1244, n_1250, n_1256 : std_logic;
  signal n_1262, n_1268, n_1274, n_1280, n_1286 : std_logic;
  signal n_1292, n_1298, n_1304, n_1310, n_1316 : std_logic;
  signal n_1322, n_1328, n_1334, n_1340, n_1346 : std_logic;
  signal n_1352, n_1358, n_1364, n_1370, n_1376 : std_logic;
  signal n_1382, n_1388, n_1394, n_1400, n_1406 : std_logic;
  signal n_1412, n_1418, n_1424, n_1430, n_1436 : std_logic;
  signal n_1442, n_1448, n_1454, n_1460, n_1466 : std_logic;
  signal n_1472, n_1478, n_1482, n_1483, n_1484 : std_logic;

begin

  counter_reg_7 : DFKCNQD1BWP7T port map(CP => clk, CN => new_counter(7), D => n_355, Q => counter(7));
  counter_reg_6 : DFKCNQD1BWP7T port map(CP => clk, CN => new_counter(6), D => n_355, Q => counter(6));
  new_counter_reg_7 : LHQD1BWP7T port map(E => n_354, D => n_352, Q => new_counter(7));
  new_counter_reg_6 : LHQD1BWP7T port map(E => n_354, D => n_353, Q => new_counter(6));
  g17264 : OAI31D0BWP7T port map(A1 => counter(6), A2 => n_299, A3 => n_305, B => n_1482, ZN => n_353);
  new_calc_buf_out_reg_3 : LHQD1BWP7T port map(E => n_351, D => n_334, Q => new_calc_buf_out(3));
  g17197 : IOA21D0BWP7T port map(A1 => n_316, A2 => counter(7), B => n_294, ZN => n_352);
  new_calc_buf_out_reg_6 : LHQD1BWP7T port map(E => n_351, D => n_340, Q => new_calc_buf_out(6));
  new_calc_buf_out_reg_7 : LHQD1BWP7T port map(E => n_351, D => n_342, Q => new_calc_buf_out(7));
  new_calc_buf_out_reg_14 : LHQD1BWP7T port map(E => n_350, D => n_346, Q => new_calc_buf_out(14));
  new_calc_buf_out_reg_15 : LHQD1BWP7T port map(E => n_350, D => n_345, Q => new_calc_buf_out(15));
  new_calc_buf_out_reg_4 : LHQD1BWP7T port map(E => n_351, D => n_333, Q => new_calc_buf_out(4));
  new_calc_buf_out_reg_5 : LHQD1BWP7T port map(E => n_351, D => n_332, Q => new_calc_buf_out(5));
  new_calc_buf_out_reg_0 : LHQD1BWP7T port map(E => n_351, D => n_319, Q => new_calc_buf_out(0));
  new_calc_buf_out_reg_1 : LHQD1BWP7T port map(E => n_351, D => n_336, Q => new_calc_buf_out(1));
  new_calc_buf_out_reg_2 : LHQD1BWP7T port map(E => n_351, D => n_335, Q => new_calc_buf_out(2));
  new_calc_buf_out_reg_9 : LHQD1BWP7T port map(E => n_350, D => n_330, Q => new_calc_buf_out(9));
  new_calc_buf_out_reg_10 : LHQD1BWP7T port map(E => n_350, D => n_328, Q => new_calc_buf_out(10));
  new_calc_buf_out_reg_11 : LHQD1BWP7T port map(E => n_350, D => n_326, Q => new_calc_buf_out(11));
  new_calc_buf_out_reg_8 : LHQD1BWP7T port map(E => n_350, D => n_331, Q => new_calc_buf_out(8));
  new_calc_buf_out_reg_12 : LHQD1BWP7T port map(E => n_350, D => n_324, Q => new_calc_buf_out(12));
  new_calc_buf_out_reg_13 : LHQD1BWP7T port map(E => n_350, D => n_322, Q => new_calc_buf_out(13));
  new_calc_buf_out_reg_18 : LHQD1BWP7T port map(E => n_350, D => n_309, Q => new_calc_buf_out(18));
  new_calc_buf_out_reg_23 : LHQD1BWP7T port map(E => n_350, D => n_307, Q => new_calc_buf_out(23));
  new_calc_buf_out_reg_16 : LHQD1BWP7T port map(E => n_350, D => n_311, Q => new_calc_buf_out(16));
  new_calc_buf_out_reg_17 : LHQD1BWP7T port map(E => n_350, D => n_310, Q => new_calc_buf_out(17));
  new_calc_buf_out_reg_22 : LHQD1BWP7T port map(E => n_350, D => n_317, Q => new_calc_buf_out(22));
  new_calc_buf_out_reg_19 : LHQD1BWP7T port map(E => n_350, D => n_308, Q => new_calc_buf_out(19));
  new_calc_buf_out_reg_20 : LHQD1BWP7T port map(E => n_350, D => n_312, Q => new_calc_buf_out(20));
  new_calc_buf_out_reg_21 : LHQD1BWP7T port map(E => n_350, D => n_315, Q => new_calc_buf_out(21));
  counter_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => new_counter(1), D => n_355, Q => counter(1));
  counter_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => new_counter(0), D => n_355, Q => counter(0));
  g17260 : MOAI22D0BWP7T port map(A1 => n_344, A2 => n_338, B1 => n_343, B2 => calc_buf_out_14_3528, ZN => n_346);
  g17259 : MOAI22D0BWP7T port map(A1 => n_344, A2 => n_341, B1 => n_343, B2 => calc_buf_out_15_3529, ZN => n_345);
  g17261 : MOAI22D0BWP7T port map(A1 => n_339, A2 => n_341, B1 => n_337, B2 => calc_buf_out_7_3521, ZN => n_342);
  new_counter_reg_5 : LHQD1BWP7T port map(E => n_354, D => n_306, Q => new_counter(5));
  new_counter_reg_3 : LHQD1BWP7T port map(E => n_354, D => n_304, Q => new_counter(3));
  g17265 : MOAI22D0BWP7T port map(A1 => n_339, A2 => n_338, B1 => n_337, B2 => calc_buf_out_6_3520, ZN => n_340);
  g17272 : MOAI22D0BWP7T port map(A1 => n_339, A2 => n_329, B1 => n_337, B2 => calc_buf_out_1_3515, ZN => n_336);
  g17273 : MOAI22D0BWP7T port map(A1 => n_339, A2 => n_327, B1 => n_337, B2 => calc_buf_out_2_3516, ZN => n_335);
  g17274 : MOAI22D0BWP7T port map(A1 => n_339, A2 => n_325, B1 => n_337, B2 => calc_buf_out_3_3517, ZN => n_334);
  g17275 : MOAI22D0BWP7T port map(A1 => n_339, A2 => n_323, B1 => n_337, B2 => calc_buf_out_4_3518, ZN => n_333);
  g17276 : MOAI22D0BWP7T port map(A1 => n_339, A2 => n_321, B1 => n_337, B2 => calc_buf_out_5_3519, ZN => n_332);
  g17277 : MOAI22D0BWP7T port map(A1 => n_344, A2 => n_318, B1 => n_343, B2 => calc_buf_out_8_3522, ZN => n_331);
  g17278 : MOAI22D0BWP7T port map(A1 => n_344, A2 => n_329, B1 => n_343, B2 => calc_buf_out_9_3523, ZN => n_330);
  g17279 : MOAI22D0BWP7T port map(A1 => n_344, A2 => n_327, B1 => n_343, B2 => calc_buf_out_10_3524, ZN => n_328);
  g17280 : MOAI22D0BWP7T port map(A1 => n_344, A2 => n_325, B1 => n_343, B2 => calc_buf_out_11_3525, ZN => n_326);
  g17281 : MOAI22D0BWP7T port map(A1 => n_344, A2 => n_323, B1 => n_343, B2 => calc_buf_out_12_3526, ZN => n_324);
  g17282 : MOAI22D0BWP7T port map(A1 => n_344, A2 => n_321, B1 => n_343, B2 => calc_buf_out_13_3527, ZN => n_322);
  g17256 : MOAI22D0BWP7T port map(A1 => n_339, A2 => n_318, B1 => n_337, B2 => calc_buf_out_0_3514, ZN => n_319);
  state_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => n_347, D => n_300, Q => state(1));
  g17258 : MOAI22D0BWP7T port map(A1 => n_314, A2 => n_338, B1 => n_313, B2 => calc_buf_out_22_3536, ZN => n_317);
  g17360 : OAI21D0BWP7T port map(A1 => n_156, A2 => counter(6), B => n_302, ZN => n_316);
  g17288 : MOAI22D0BWP7T port map(A1 => n_314, A2 => n_321, B1 => n_313, B2 => calc_buf_out_21_3535, ZN => n_315);
  g17287 : MOAI22D0BWP7T port map(A1 => n_314, A2 => n_323, B1 => n_313, B2 => calc_buf_out_20_3534, ZN => n_312);
  g17283 : MOAI22D0BWP7T port map(A1 => n_314, A2 => n_318, B1 => n_313, B2 => calc_buf_out_16_3530, ZN => n_311);
  g17284 : MOAI22D0BWP7T port map(A1 => n_314, A2 => n_329, B1 => n_313, B2 => calc_buf_out_17_3531, ZN => n_310);
  g17285 : MOAI22D0BWP7T port map(A1 => n_314, A2 => n_327, B1 => n_313, B2 => calc_buf_out_18_3532, ZN => n_309);
  g17286 : MOAI22D0BWP7T port map(A1 => n_314, A2 => n_325, B1 => n_313, B2 => calc_buf_out_19_3533, ZN => n_308);
  state_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => n_347, D => n_288, Q => state(0));
  g17257 : MOAI22D0BWP7T port map(A1 => n_314, A2 => n_341, B1 => n_313, B2 => calc_buf_out_23_3537, ZN => n_307);
  g17326 : MOAI22D0BWP7T port map(A1 => n_305, A2 => counter(5), B1 => n_298, B2 => counter(5), ZN => n_306);
  new_counter_reg_1 : LHQD1BWP7T port map(E => n_354, D => n_291, Q => new_counter(1));
  g17359 : AO21D0BWP7T port map(A1 => n_157, A2 => counter(3), B => n_75, Z => n_304);
  new_counter_reg_0 : LHQD1BWP7T port map(E => n_354, D => n_293, Q => new_counter(0));
  new_counter_reg_2 : LHQD1BWP7T port map(E => n_354, D => n_289, Q => new_counter(2));
  new_counter_reg_4 : LHQD1BWP7T port map(E => n_354, D => n_287, Q => new_counter(4));
  state_reg_3 : DFQD1BWP7T port map(CP => clk, D => n_281, Q => state(3));
  new_framebuffer_buf_reg_10 : LHQD1BWP7T port map(E => n_301, D => n_280, Q => new_framebuffer_buf(10));
  new_framebuffer_buf_reg_14 : LHQD1BWP7T port map(E => n_301, D => n_279, Q => new_framebuffer_buf(14));
  new_framebuffer_buf_reg_15 : LHQD1BWP7T port map(E => n_301, D => n_278, Q => new_framebuffer_buf(15));
  new_framebuffer_buf_reg_8 : LHQD1BWP7T port map(E => n_301, D => n_282, Q => new_framebuffer_buf(8));
  new_framebuffer_buf_reg_12 : LHQD1BWP7T port map(E => n_301, D => n_277, Q => new_framebuffer_buf(12));
  new_framebuffer_buf_reg_9 : LHQD1BWP7T port map(E => n_301, D => n_283, Q => new_framebuffer_buf(9));
  new_framebuffer_buf_reg_11 : LHQD1BWP7T port map(E => n_301, D => n_296, Q => new_framebuffer_buf(11));
  new_framebuffer_buf_reg_13 : LHQD1BWP7T port map(E => n_301, D => n_284, Q => new_framebuffer_buf(13));
  new_framebuffer_buf_reg_100 : LHQD1BWP7T port map(E => n_301, D => n_255, Q => new_framebuffer_buf(100));
  new_framebuffer_buf_reg_101 : LHQD1BWP7T port map(E => n_301, D => n_254, Q => new_framebuffer_buf(101));
  new_framebuffer_buf_reg_104 : LHQD1BWP7T port map(E => n_301, D => n_253, Q => new_framebuffer_buf(104));
  new_framebuffer_buf_reg_105 : LHQD1BWP7T port map(E => n_301, D => n_252, Q => new_framebuffer_buf(105));
  new_framebuffer_buf_reg_106 : LHQD1BWP7T port map(E => n_301, D => n_251, Q => new_framebuffer_buf(106));
  new_framebuffer_buf_reg_107 : LHQD1BWP7T port map(E => n_301, D => n_260, Q => new_framebuffer_buf(107));
  new_framebuffer_buf_reg_108 : LHQD1BWP7T port map(E => n_301, D => n_248, Q => new_framebuffer_buf(108));
  new_framebuffer_buf_reg_109 : LHQD1BWP7T port map(E => n_301, D => n_247, Q => new_framebuffer_buf(109));
  new_framebuffer_buf_reg_112 : LHQD1BWP7T port map(E => n_301, D => n_245, Q => new_framebuffer_buf(112));
  new_framebuffer_buf_reg_113 : LHQD1BWP7T port map(E => n_301, D => n_244, Q => new_framebuffer_buf(113));
  new_framebuffer_buf_reg_114 : LHQD1BWP7T port map(E => n_301, D => n_242, Q => new_framebuffer_buf(114));
  new_framebuffer_buf_reg_116 : LHQD1BWP7T port map(E => n_301, D => n_241, Q => new_framebuffer_buf(116));
  new_framebuffer_buf_reg_117 : LHQD1BWP7T port map(E => n_301, D => n_240, Q => new_framebuffer_buf(117));
  new_framebuffer_buf_reg_120 : LHQD1BWP7T port map(E => n_301, D => n_270, Q => new_framebuffer_buf(120));
  new_framebuffer_buf_reg_122 : LHQD1BWP7T port map(E => n_301, D => n_274, Q => new_framebuffer_buf(122));
  new_framebuffer_buf_reg_123 : LHQD1BWP7T port map(E => n_301, D => n_272, Q => new_framebuffer_buf(123));
  new_framebuffer_buf_reg_124 : LHQD1BWP7T port map(E => n_301, D => n_142, Q => new_framebuffer_buf(124));
  new_framebuffer_buf_reg_125 : LHQD1BWP7T port map(E => n_301, D => n_271, Q => new_framebuffer_buf(125));
  new_framebuffer_buf_reg_56 : LHQD1BWP7T port map(E => n_301, D => n_209, Q => new_framebuffer_buf(56));
  new_framebuffer_buf_reg_38 : LHQD1BWP7T port map(E => n_301, D => n_169, Q => new_framebuffer_buf(38));
  new_framebuffer_buf_reg_39 : LHQD1BWP7T port map(E => n_301, D => n_168, Q => new_framebuffer_buf(39));
  new_framebuffer_buf_reg_46 : LHQD1BWP7T port map(E => n_301, D => n_191, Q => new_framebuffer_buf(46));
  new_framebuffer_buf_reg_47 : LHQD1BWP7T port map(E => n_301, D => n_190, Q => new_framebuffer_buf(47));
  new_framebuffer_buf_reg_54 : LHQD1BWP7T port map(E => n_301, D => n_189, Q => new_framebuffer_buf(54));
  new_framebuffer_buf_reg_55 : LHQD1BWP7T port map(E => n_301, D => n_187, Q => new_framebuffer_buf(55));
  new_framebuffer_buf_reg_62 : LHQD1BWP7T port map(E => n_301, D => n_218, Q => new_framebuffer_buf(62));
  new_framebuffer_buf_reg_63 : LHQD1BWP7T port map(E => n_301, D => n_216, Q => new_framebuffer_buf(63));
  new_framebuffer_buf_reg_70 : LHQD1BWP7T port map(E => n_301, D => n_172, Q => new_framebuffer_buf(70));
  new_framebuffer_buf_reg_71 : LHQD1BWP7T port map(E => n_301, D => n_170, Q => new_framebuffer_buf(71));
  new_framebuffer_buf_reg_78 : LHQD1BWP7T port map(E => n_301, D => n_215, Q => new_framebuffer_buf(78));
  new_framebuffer_buf_reg_79 : LHQD1BWP7T port map(E => n_301, D => n_213, Q => new_framebuffer_buf(79));
  new_framebuffer_buf_reg_86 : LHQD1BWP7T port map(E => n_301, D => n_212, Q => new_framebuffer_buf(86));
  new_framebuffer_buf_reg_87 : LHQD1BWP7T port map(E => n_301, D => n_210, Q => new_framebuffer_buf(87));
  new_framebuffer_buf_reg_94 : LHQD1BWP7T port map(E => n_301, D => n_230, Q => new_framebuffer_buf(94));
  new_framebuffer_buf_reg_95 : LHQD1BWP7T port map(E => n_301, D => n_228, Q => new_framebuffer_buf(95));
  new_framebuffer_buf_reg_32 : LHQD1BWP7T port map(E => n_301, D => n_161, Q => new_framebuffer_buf(32));
  new_framebuffer_buf_reg_33 : LHQD1BWP7T port map(E => n_301, D => n_160, Q => new_framebuffer_buf(33));
  new_framebuffer_buf_reg_34 : LHQD1BWP7T port map(E => n_301, D => n_159, Q => new_framebuffer_buf(34));
  new_framebuffer_buf_reg_35 : LHQD1BWP7T port map(E => n_301, D => n_243, Q => new_framebuffer_buf(35));
  new_framebuffer_buf_reg_36 : LHQD1BWP7T port map(E => n_301, D => n_246, Q => new_framebuffer_buf(36));
  new_framebuffer_buf_reg_37 : LHQD1BWP7T port map(E => n_301, D => n_250, Q => new_framebuffer_buf(37));
  new_framebuffer_buf_reg_40 : LHQD1BWP7T port map(E => n_301, D => n_220, Q => new_framebuffer_buf(40));
  new_framebuffer_buf_reg_41 : LHQD1BWP7T port map(E => n_301, D => n_222, Q => new_framebuffer_buf(41));
  new_framebuffer_buf_reg_42 : LHQD1BWP7T port map(E => n_301, D => n_153, Q => new_framebuffer_buf(42));
  new_framebuffer_buf_reg_43 : LHQD1BWP7T port map(E => n_301, D => n_183, Q => new_framebuffer_buf(43));
  new_framebuffer_buf_reg_44 : LHQD1BWP7T port map(E => n_301, D => n_182, Q => new_framebuffer_buf(44));
  new_framebuffer_buf_reg_45 : LHQD1BWP7T port map(E => n_301, D => n_179, Q => new_framebuffer_buf(45));
  g17209 : ND4D0BWP7T port map(A1 => n_125, A2 => n_73, A3 => n_48, A4 => n_28, ZN => n_300);
  new_framebuffer_buf_reg_48 : LHQD1BWP7T port map(E => n_301, D => n_178, Q => new_framebuffer_buf(48));
  new_framebuffer_buf_reg_49 : LHQD1BWP7T port map(E => n_301, D => n_177, Q => new_framebuffer_buf(49));
  new_framebuffer_buf_reg_50 : LHQD1BWP7T port map(E => n_301, D => n_176, Q => new_framebuffer_buf(50));
  new_framebuffer_buf_reg_51 : LHQD1BWP7T port map(E => n_301, D => n_175, Q => new_framebuffer_buf(51));
  new_framebuffer_buf_reg_52 : LHQD1BWP7T port map(E => n_301, D => n_174, Q => new_framebuffer_buf(52));
  new_framebuffer_buf_reg_53 : LHQD1BWP7T port map(E => n_301, D => n_173, Q => new_framebuffer_buf(53));
  new_framebuffer_buf_reg_58 : LHQD1BWP7T port map(E => n_301, D => n_207, Q => new_framebuffer_buf(58));
  new_framebuffer_buf_reg_59 : LHQD1BWP7T port map(E => n_301, D => n_206, Q => new_framebuffer_buf(59));
  new_framebuffer_buf_reg_60 : LHQD1BWP7T port map(E => n_301, D => n_205, Q => new_framebuffer_buf(60));
  new_framebuffer_buf_reg_61 : LHQD1BWP7T port map(E => n_301, D => n_204, Q => new_framebuffer_buf(61));
  new_framebuffer_buf_reg_64 : LHQD1BWP7T port map(E => n_301, D => n_167, Q => new_framebuffer_buf(64));
  new_framebuffer_buf_reg_65 : LHQD1BWP7T port map(E => n_301, D => n_166, Q => new_framebuffer_buf(65));
  new_framebuffer_buf_reg_66 : LHQD1BWP7T port map(E => n_301, D => n_165, Q => new_framebuffer_buf(66));
  g17525 : AOI21D0BWP7T port map(A1 => n_122, A2 => n_299, B => n_298, ZN => n_302);
  new_framebuffer_buf_reg_67 : LHQD1BWP7T port map(E => n_301, D => n_164, Q => new_framebuffer_buf(67));
  new_framebuffer_buf_reg_99 : LHQD1BWP7T port map(E => n_301, D => n_256, Q => new_framebuffer_buf(99));
  new_framebuffer_buf_reg_68 : LHQD1BWP7T port map(E => n_301, D => n_163, Q => new_framebuffer_buf(68));
  new_framebuffer_buf_reg_69 : LHQD1BWP7T port map(E => n_301, D => n_162, Q => new_framebuffer_buf(69));
  new_framebuffer_buf_reg_72 : LHQD1BWP7T port map(E => n_301, D => n_203, Q => new_framebuffer_buf(72));
  new_framebuffer_buf_reg_98 : LHQD1BWP7T port map(E => n_301, D => n_257, Q => new_framebuffer_buf(98));
  new_framebuffer_buf_reg_73 : LHQD1BWP7T port map(E => n_301, D => n_202, Q => new_framebuffer_buf(73));
  new_framebuffer_buf_reg_74 : LHQD1BWP7T port map(E => n_301, D => n_201, Q => new_framebuffer_buf(74));
  new_framebuffer_buf_reg_75 : LHQD1BWP7T port map(E => n_301, D => n_200, Q => new_framebuffer_buf(75));
  new_framebuffer_buf_reg_76 : LHQD1BWP7T port map(E => n_301, D => n_199, Q => new_framebuffer_buf(76));
  new_framebuffer_buf_reg_77 : LHQD1BWP7T port map(E => n_301, D => n_198, Q => new_framebuffer_buf(77));
  new_framebuffer_buf_reg_80 : LHQD1BWP7T port map(E => n_301, D => n_197, Q => new_framebuffer_buf(80));
  new_framebuffer_buf_reg_81 : LHQD1BWP7T port map(E => n_301, D => n_196, Q => new_framebuffer_buf(81));
  new_framebuffer_buf_reg_82 : LHQD1BWP7T port map(E => n_301, D => n_195, Q => new_framebuffer_buf(82));
  new_framebuffer_buf_reg_83 : LHQD1BWP7T port map(E => n_301, D => n_194, Q => new_framebuffer_buf(83));
  new_framebuffer_buf_reg_84 : LHQD1BWP7T port map(E => n_301, D => n_193, Q => new_framebuffer_buf(84));
  new_framebuffer_buf_reg_85 : LHQD1BWP7T port map(E => n_301, D => n_192, Q => new_framebuffer_buf(85));
  new_framebuffer_buf_reg_88 : LHQD1BWP7T port map(E => n_301, D => n_227, Q => new_framebuffer_buf(88));
  new_framebuffer_buf_reg_89 : LHQD1BWP7T port map(E => n_301, D => n_226, Q => new_framebuffer_buf(89));
  new_framebuffer_buf_reg_90 : LHQD1BWP7T port map(E => n_301, D => n_225, Q => new_framebuffer_buf(90));
  new_framebuffer_buf_reg_91 : LHQD1BWP7T port map(E => n_301, D => n_224, Q => new_framebuffer_buf(91));
  new_framebuffer_buf_reg_92 : LHQD1BWP7T port map(E => n_301, D => n_223, Q => new_framebuffer_buf(92));
  new_framebuffer_buf_reg_93 : LHQD1BWP7T port map(E => n_301, D => n_219, Q => new_framebuffer_buf(93));
  new_framebuffer_buf_reg_57 : LHQD1BWP7T port map(E => n_301, D => n_208, Q => new_framebuffer_buf(57));
  new_framebuffer_buf_reg_30 : LHQD1BWP7T port map(E => n_301, D => n_181, Q => new_framebuffer_buf(30));
  new_framebuffer_buf_reg_31 : LHQD1BWP7T port map(E => n_301, D => n_158, Q => new_framebuffer_buf(31));
  new_framebuffer_buf_reg_25 : LHQD1BWP7T port map(E => n_301, D => n_151, Q => new_framebuffer_buf(25));
  new_framebuffer_buf_reg_26 : LHQD1BWP7T port map(E => n_301, D => n_150, Q => new_framebuffer_buf(26));
  new_framebuffer_buf_reg_27 : LHQD1BWP7T port map(E => n_301, D => n_149, Q => new_framebuffer_buf(27));
  new_framebuffer_buf_reg_28 : LHQD1BWP7T port map(E => n_301, D => n_148, Q => new_framebuffer_buf(28));
  new_framebuffer_buf_reg_29 : LHQD1BWP7T port map(E => n_301, D => n_147, Q => new_framebuffer_buf(29));
  new_framebuffer_buf_reg_24 : LHQD1BWP7T port map(E => n_301, D => n_152, Q => new_framebuffer_buf(24));
  new_framebuffer_buf_reg_22 : LHQD1BWP7T port map(E => n_301, D => n_146, Q => new_framebuffer_buf(22));
  new_framebuffer_buf_reg_23 : LHQD1BWP7T port map(E => n_301, D => n_144, Q => new_framebuffer_buf(23));
  new_framebuffer_buf_reg_115 : LHQD1BWP7T port map(E => n_301, D => n_259, Q => new_framebuffer_buf(115));
  new_framebuffer_buf_reg_16 : LHQD1BWP7T port map(E => n_301, D => n_141, Q => new_framebuffer_buf(16));
  new_framebuffer_buf_reg_17 : LHQD1BWP7T port map(E => n_301, D => n_140, Q => new_framebuffer_buf(17));
  new_framebuffer_buf_reg_18 : LHQD1BWP7T port map(E => n_301, D => n_139, Q => new_framebuffer_buf(18));
  new_framebuffer_buf_reg_19 : LHQD1BWP7T port map(E => n_301, D => n_138, Q => new_framebuffer_buf(19));
  new_framebuffer_buf_reg_20 : LHQD1BWP7T port map(E => n_301, D => n_137, Q => new_framebuffer_buf(20));
  new_framebuffer_buf_reg_21 : LHQD1BWP7T port map(E => n_301, D => n_136, Q => new_framebuffer_buf(21));
  new_framebuffer_buf_reg_6 : LHQD1BWP7T port map(E => n_301, D => n_135, Q => new_framebuffer_buf(6));
  new_framebuffer_buf_reg_7 : LHQD1BWP7T port map(E => n_301, D => n_133, Q => new_framebuffer_buf(7));
  new_framebuffer_buf_reg_0 : LHQD1BWP7T port map(E => n_301, D => n_132, Q => new_framebuffer_buf(0));
  new_framebuffer_buf_reg_1 : LHQD1BWP7T port map(E => n_301, D => n_131, Q => new_framebuffer_buf(1));
  new_framebuffer_buf_reg_2 : LHQD1BWP7T port map(E => n_301, D => n_130, Q => new_framebuffer_buf(2));
  new_framebuffer_buf_reg_3 : LHQD1BWP7T port map(E => n_301, D => n_129, Q => new_framebuffer_buf(3));
  new_framebuffer_buf_reg_4 : LHQD1BWP7T port map(E => n_301, D => n_128, Q => new_framebuffer_buf(4));
  new_framebuffer_buf_reg_5 : LHQD1BWP7T port map(E => n_301, D => n_127, Q => new_framebuffer_buf(5));
  new_framebuffer_buf_reg_127 : LHQD1BWP7T port map(E => n_301, D => n_154, Q => new_framebuffer_buf(127));
  new_framebuffer_buf_reg_118 : LHQD1BWP7T port map(E => n_301, D => n_263, Q => new_framebuffer_buf(118));
  new_framebuffer_buf_reg_102 : LHQD1BWP7T port map(E => n_301, D => n_267, Q => new_framebuffer_buf(102));
  new_framebuffer_buf_reg_103 : LHQD1BWP7T port map(E => n_301, D => n_265, Q => new_framebuffer_buf(103));
  new_framebuffer_buf_reg_110 : LHQD1BWP7T port map(E => n_301, D => n_269, Q => new_framebuffer_buf(110));
  new_framebuffer_buf_reg_111 : LHQD1BWP7T port map(E => n_301, D => n_264, Q => new_framebuffer_buf(111));
  new_framebuffer_buf_reg_119 : LHQD1BWP7T port map(E => n_301, D => n_261, Q => new_framebuffer_buf(119));
  new_framebuffer_buf_reg_126 : LHQD1BWP7T port map(E => n_301, D => n_143, Q => new_framebuffer_buf(126));
  new_framebuffer_buf_reg_121 : LHQD1BWP7T port map(E => n_301, D => n_231, Q => new_framebuffer_buf(121));
  new_framebuffer_buf_reg_96 : LHQD1BWP7T port map(E => n_301, D => n_239, Q => new_framebuffer_buf(96));
  new_framebuffer_buf_reg_97 : LHQD1BWP7T port map(E => n_301, D => n_258, Q => new_framebuffer_buf(97));
  g17528 : OAI21D0BWP7T port map(A1 => n_285, A2 => n_297, B => n_286, ZN => n_343);
  g17527 : OAI221D0BWP7T port map(A1 => n_65, A2 => n_292, B1 => n_297, B2 => n_186, C => n_116, ZN => n_337);
  g17604 : MOAI22D0BWP7T port map(A1 => n_1483, A2 => n_325, B1 => n_1483, B2 => framebuffer_buf_11_3549, ZN => n_296);
  g17456 : IIND4D0BWP7T port map(A1 => n_305, A2 => counter(7), B1 => counter(6), B2 => counter(5), ZN => n_294);
  g17457 : OAI221D0BWP7T port map(A1 => n_66, A2 => n_292, B1 => counter(0), B2 => n_290, C => n_115, ZN => n_293);
  g17462 : OAI21D0BWP7T port map(A1 => n_290, A2 => n_93, B => n_123, ZN => n_291);
  g17463 : OAI32D0BWP7T port map(A1 => counter(2), A2 => n_95, A3 => n_290, B1 => n_74, B2 => n_155, ZN => n_289);
  g17196 : IND4D0BWP7T port map(A1 => n_104, B1 => n_72, B2 => n_51, B3 => n_118, ZN => n_288);
  g17454 : OAI22D0BWP7T port map(A1 => n_126, A2 => n_13, B1 => n_94, B2 => counter(4), ZN => n_287);
  g17526 : OAI21D0BWP7T port map(A1 => n_184, A2 => n_297, B => n_286, ZN => n_313);
  g17667 : ND2D0BWP7T port map(A1 => n_285, A2 => n_185, ZN => n_344);
  g17581 : MOAI22D0BWP7T port map(A1 => n_1483, A2 => n_321, B1 => n_1483, B2 => framebuffer_buf_13_3551, ZN => n_284);
  g17538 : MOAI22D0BWP7T port map(A1 => n_1483, A2 => n_329, B1 => n_1483, B2 => framebuffer_buf_9_3547, ZN => n_283);
  g17539 : MOAI22D0BWP7T port map(A1 => n_1483, A2 => n_318, B1 => n_1483, B2 => framebuffer_buf_8_3546, ZN => n_282);
  g17223 : ND4D0BWP7T port map(A1 => n_106, A2 => n_20, A3 => n_276, A4 => n_355, ZN => n_281);
  g17535 : MOAI22D0BWP7T port map(A1 => n_1483, A2 => n_327, B1 => n_1483, B2 => framebuffer_buf_10_3548, ZN => n_280);
  g17572 : MOAI22D0BWP7T port map(A1 => n_1483, A2 => n_338, B1 => n_1483, B2 => framebuffer_buf_14_3552, ZN => n_279);
  g17573 : MOAI22D0BWP7T port map(A1 => n_1483, A2 => n_341, B1 => n_1483, B2 => framebuffer_buf_15_3553, ZN => n_278);
  g17580 : MOAI22D0BWP7T port map(A1 => n_1483, A2 => n_323, B1 => n_1483, B2 => framebuffer_buf_12_3550, ZN => n_277);
  g17362 : ND3D0BWP7T port map(A1 => n_286, A2 => n_297, A3 => n_276, ZN => n_350);
  g17646 : CKND4BWP7T port map(I => n_362, ZN => sqi_data_out(2));
  g17600 : MOAI22D0BWP7T port map(A1 => n_273, A2 => n_327, B1 => n_273, B2 => framebuffer_buf_122_3660, ZN => n_274);
  g17601 : MOAI22D0BWP7T port map(A1 => n_273, A2 => n_325, B1 => n_273, B2 => framebuffer_buf_123_3661, ZN => n_272);
  g17602 : MOAI22D0BWP7T port map(A1 => n_273, A2 => n_321, B1 => n_273, B2 => framebuffer_buf_125_3663, ZN => n_271);
  g17603 : MOAI22D0BWP7T port map(A1 => n_273, A2 => n_318, B1 => n_273, B2 => framebuffer_buf_120_3658, ZN => n_270);
  g17605 : MOAI22D0BWP7T port map(A1 => n_268, A2 => n_338, B1 => n_268, B2 => framebuffer_buf_110_3648, ZN => n_269);
  g17606 : MOAI22D0BWP7T port map(A1 => n_266, A2 => n_338, B1 => n_266, B2 => framebuffer_buf_102_3640, ZN => n_267);
  g17607 : MOAI22D0BWP7T port map(A1 => n_266, A2 => n_341, B1 => n_266, B2 => framebuffer_buf_103_3641, ZN => n_265);
  g17608 : MOAI22D0BWP7T port map(A1 => n_268, A2 => n_341, B1 => n_268, B2 => framebuffer_buf_111_3649, ZN => n_264);
  g17609 : MOAI22D0BWP7T port map(A1 => n_262, A2 => n_338, B1 => n_262, B2 => framebuffer_buf_118_3656, ZN => n_263);
  g17610 : MOAI22D0BWP7T port map(A1 => n_262, A2 => n_341, B1 => n_262, B2 => framebuffer_buf_119_3657, ZN => n_261);
  g17611 : MOAI22D0BWP7T port map(A1 => n_268, A2 => n_325, B1 => n_268, B2 => framebuffer_buf_107_3645, ZN => n_260);
  g17612 : MOAI22D0BWP7T port map(A1 => n_262, A2 => n_325, B1 => n_262, B2 => framebuffer_buf_115_3653, ZN => n_259);
  g17613 : MOAI22D0BWP7T port map(A1 => n_266, A2 => n_329, B1 => n_266, B2 => framebuffer_buf_97_3635, ZN => n_258);
  g17614 : MOAI22D0BWP7T port map(A1 => n_266, A2 => n_327, B1 => n_266, B2 => framebuffer_buf_98_3636, ZN => n_257);
  g17615 : MOAI22D0BWP7T port map(A1 => n_266, A2 => n_325, B1 => n_266, B2 => framebuffer_buf_99_3637, ZN => n_256);
  g17616 : MOAI22D0BWP7T port map(A1 => n_266, A2 => n_323, B1 => n_266, B2 => framebuffer_buf_100_3638, ZN => n_255);
  g17617 : MOAI22D0BWP7T port map(A1 => n_266, A2 => n_321, B1 => n_266, B2 => framebuffer_buf_101_3639, ZN => n_254);
  g17618 : MOAI22D0BWP7T port map(A1 => n_268, A2 => n_318, B1 => n_268, B2 => framebuffer_buf_104_3642, ZN => n_253);
  g17619 : MOAI22D0BWP7T port map(A1 => n_268, A2 => n_329, B1 => n_268, B2 => framebuffer_buf_105_3643, ZN => n_252);
  g17620 : MOAI22D0BWP7T port map(A1 => n_268, A2 => n_327, B1 => n_268, B2 => framebuffer_buf_106_3644, ZN => n_251);
  g17458 : MOAI22D0BWP7T port map(A1 => n_249, A2 => n_321, B1 => n_249, B2 => framebuffer_buf_37_3575, ZN => n_250);
  g17621 : MOAI22D0BWP7T port map(A1 => n_268, A2 => n_323, B1 => n_268, B2 => framebuffer_buf_108_3646, ZN => n_248);
  g17622 : MOAI22D0BWP7T port map(A1 => n_268, A2 => n_321, B1 => n_268, B2 => framebuffer_buf_109_3647, ZN => n_247);
  g17459 : MOAI22D0BWP7T port map(A1 => n_249, A2 => n_323, B1 => n_249, B2 => framebuffer_buf_36_3574, ZN => n_246);
  g17623 : MOAI22D0BWP7T port map(A1 => n_262, A2 => n_318, B1 => n_262, B2 => framebuffer_buf_112_3650, ZN => n_245);
  g17624 : MOAI22D0BWP7T port map(A1 => n_262, A2 => n_329, B1 => n_262, B2 => framebuffer_buf_113_3651, ZN => n_244);
  g17460 : MOAI22D0BWP7T port map(A1 => n_249, A2 => n_325, B1 => n_249, B2 => framebuffer_buf_35_3573, ZN => n_243);
  g17625 : MOAI22D0BWP7T port map(A1 => n_262, A2 => n_327, B1 => n_262, B2 => framebuffer_buf_114_3652, ZN => n_242);
  g17626 : MOAI22D0BWP7T port map(A1 => n_262, A2 => n_323, B1 => n_262, B2 => framebuffer_buf_116_3654, ZN => n_241);
  g17627 : MOAI22D0BWP7T port map(A1 => n_262, A2 => n_321, B1 => n_262, B2 => framebuffer_buf_117_3655, ZN => n_240);
  g17628 : MOAI22D0BWP7T port map(A1 => n_266, A2 => n_318, B1 => n_266, B2 => framebuffer_buf_96_3634, ZN => n_239);
  new_framebuffer_buf_reg_152 : LHQD1BWP7T port map(E => n_301, D => n_109, Q => new_framebuffer_buf(152));
  g17631 : CKND4BWP7T port map(I => n_369, ZN => sqi_data_out(6));
  g17634 : CKND4BWP7T port map(I => n_368, ZN => sqi_data_out(7));
  g17636 : CKND4BWP7T port map(I => n_367, ZN => sqi_data_out(0));
  g17638 : CKND4BWP7T port map(I => n_366, ZN => sqi_data_out(5));
  g17640 : CKND4BWP7T port map(I => n_365, ZN => sqi_data_out(1));
  g17642 : CKND4BWP7T port map(I => n_364, ZN => sqi_data_out(4));
  g17644 : CKND4BWP7T port map(I => n_363, ZN => sqi_data_out(3));
  g17599 : MOAI22D0BWP7T port map(A1 => n_273, A2 => n_329, B1 => n_273, B2 => framebuffer_buf_121_3659, ZN => n_231);
  g17464 : MOAI22D0BWP7T port map(A1 => n_229, A2 => n_338, B1 => n_229, B2 => framebuffer_buf_94_3632, ZN => n_230);
  g17465 : MOAI22D0BWP7T port map(A1 => n_229, A2 => n_341, B1 => n_229, B2 => framebuffer_buf_95_3633, ZN => n_228);
  g17466 : MOAI22D0BWP7T port map(A1 => n_229, A2 => n_318, B1 => n_229, B2 => framebuffer_buf_88_3626, ZN => n_227);
  g17467 : MOAI22D0BWP7T port map(A1 => n_229, A2 => n_329, B1 => n_229, B2 => framebuffer_buf_89_3627, ZN => n_226);
  g17468 : MOAI22D0BWP7T port map(A1 => n_229, A2 => n_327, B1 => n_229, B2 => framebuffer_buf_90_3628, ZN => n_225);
  g17469 : MOAI22D0BWP7T port map(A1 => n_229, A2 => n_325, B1 => n_229, B2 => framebuffer_buf_91_3629, ZN => n_224);
  g17470 : MOAI22D0BWP7T port map(A1 => n_229, A2 => n_323, B1 => n_229, B2 => framebuffer_buf_92_3630, ZN => n_223);
  g17501 : MOAI22D0BWP7T port map(A1 => n_221, A2 => n_329, B1 => n_221, B2 => framebuffer_buf_41_3579, ZN => n_222);
  g17500 : MOAI22D0BWP7T port map(A1 => n_221, A2 => n_318, B1 => n_221, B2 => framebuffer_buf_40_3578, ZN => n_220);
  g17471 : MOAI22D0BWP7T port map(A1 => n_229, A2 => n_321, B1 => n_229, B2 => framebuffer_buf_93_3631, ZN => n_219);
  g17472 : MOAI22D0BWP7T port map(A1 => n_217, A2 => n_338, B1 => n_217, B2 => framebuffer_buf_62_3600, ZN => n_218);
  g17473 : MOAI22D0BWP7T port map(A1 => n_217, A2 => n_341, B1 => n_217, B2 => framebuffer_buf_63_3601, ZN => n_216);
  g17474 : MOAI22D0BWP7T port map(A1 => n_214, A2 => n_338, B1 => n_214, B2 => framebuffer_buf_78_3616, ZN => n_215);
  g17475 : MOAI22D0BWP7T port map(A1 => n_214, A2 => n_341, B1 => n_214, B2 => framebuffer_buf_79_3617, ZN => n_213);
  g17476 : MOAI22D0BWP7T port map(A1 => n_211, A2 => n_338, B1 => n_211, B2 => framebuffer_buf_86_3624, ZN => n_212);
  g17477 : MOAI22D0BWP7T port map(A1 => n_211, A2 => n_341, B1 => n_211, B2 => framebuffer_buf_87_3625, ZN => n_210);
  g17478 : MOAI22D0BWP7T port map(A1 => n_217, A2 => n_318, B1 => n_217, B2 => framebuffer_buf_56_3594, ZN => n_209);
  g17479 : MOAI22D0BWP7T port map(A1 => n_217, A2 => n_329, B1 => n_217, B2 => framebuffer_buf_57_3595, ZN => n_208);
  g17480 : MOAI22D0BWP7T port map(A1 => n_217, A2 => n_327, B1 => n_217, B2 => framebuffer_buf_58_3596, ZN => n_207);
  g17481 : MOAI22D0BWP7T port map(A1 => n_217, A2 => n_325, B1 => n_217, B2 => framebuffer_buf_59_3597, ZN => n_206);
  g17482 : MOAI22D0BWP7T port map(A1 => n_217, A2 => n_323, B1 => n_217, B2 => framebuffer_buf_60_3598, ZN => n_205);
  g17483 : MOAI22D0BWP7T port map(A1 => n_217, A2 => n_321, B1 => n_217, B2 => framebuffer_buf_61_3599, ZN => n_204);
  g17484 : MOAI22D0BWP7T port map(A1 => n_214, A2 => n_318, B1 => n_214, B2 => framebuffer_buf_72_3610, ZN => n_203);
  g17485 : MOAI22D0BWP7T port map(A1 => n_214, A2 => n_329, B1 => n_214, B2 => framebuffer_buf_73_3611, ZN => n_202);
  g17486 : MOAI22D0BWP7T port map(A1 => n_214, A2 => n_327, B1 => n_214, B2 => framebuffer_buf_74_3612, ZN => n_201);
  g17487 : MOAI22D0BWP7T port map(A1 => n_214, A2 => n_325, B1 => n_214, B2 => framebuffer_buf_75_3613, ZN => n_200);
  g17488 : MOAI22D0BWP7T port map(A1 => n_214, A2 => n_323, B1 => n_214, B2 => framebuffer_buf_76_3614, ZN => n_199);
  g17489 : MOAI22D0BWP7T port map(A1 => n_214, A2 => n_321, B1 => n_214, B2 => framebuffer_buf_77_3615, ZN => n_198);
  g17490 : MOAI22D0BWP7T port map(A1 => n_211, A2 => n_318, B1 => n_211, B2 => framebuffer_buf_80_3618, ZN => n_197);
  g17491 : MOAI22D0BWP7T port map(A1 => n_211, A2 => n_329, B1 => n_211, B2 => framebuffer_buf_81_3619, ZN => n_196);
  g17492 : MOAI22D0BWP7T port map(A1 => n_211, A2 => n_327, B1 => n_211, B2 => framebuffer_buf_82_3620, ZN => n_195);
  g17493 : MOAI22D0BWP7T port map(A1 => n_211, A2 => n_325, B1 => n_211, B2 => framebuffer_buf_83_3621, ZN => n_194);
  g17494 : MOAI22D0BWP7T port map(A1 => n_211, A2 => n_323, B1 => n_211, B2 => framebuffer_buf_84_3622, ZN => n_193);
  g17495 : MOAI22D0BWP7T port map(A1 => n_211, A2 => n_321, B1 => n_211, B2 => framebuffer_buf_85_3623, ZN => n_192);
  g17496 : MOAI22D0BWP7T port map(A1 => n_221, A2 => n_338, B1 => n_221, B2 => framebuffer_buf_46_3584, ZN => n_191);
  g17497 : MOAI22D0BWP7T port map(A1 => n_221, A2 => n_341, B1 => n_221, B2 => framebuffer_buf_47_3585, ZN => n_190);
  g17498 : MOAI22D0BWP7T port map(A1 => n_188, A2 => n_338, B1 => n_188, B2 => framebuffer_buf_54_3592, ZN => n_189);
  g17499 : MOAI22D0BWP7T port map(A1 => n_188, A2 => n_341, B1 => n_188, B2 => framebuffer_buf_55_3593, ZN => n_187);
  g17668 : ND2D0BWP7T port map(A1 => n_186, A2 => n_185, ZN => n_339);
  g17666 : ND2D0BWP7T port map(A1 => n_184, A2 => n_185, ZN => n_314);
  new_framebuffer_buf_reg_141 : LHQD1BWP7T port map(E => n_301, D => n_82, Q => new_framebuffer_buf(141));
  g17503 : MOAI22D0BWP7T port map(A1 => n_221, A2 => n_325, B1 => n_221, B2 => framebuffer_buf_43_3581, ZN => n_183);
  g17504 : MOAI22D0BWP7T port map(A1 => n_221, A2 => n_323, B1 => n_221, B2 => framebuffer_buf_44_3582, ZN => n_182);
  g17558 : MOAI22D0BWP7T port map(A1 => n_180, A2 => n_338, B1 => n_180, B2 => framebuffer_buf_30_3568, ZN => n_181);
  g17505 : MOAI22D0BWP7T port map(A1 => n_221, A2 => n_321, B1 => n_221, B2 => framebuffer_buf_45_3583, ZN => n_179);
  g17506 : MOAI22D0BWP7T port map(A1 => n_188, A2 => n_318, B1 => n_188, B2 => framebuffer_buf_48_3586, ZN => n_178);
  g17507 : MOAI22D0BWP7T port map(A1 => n_188, A2 => n_329, B1 => n_188, B2 => framebuffer_buf_49_3587, ZN => n_177);
  g17508 : MOAI22D0BWP7T port map(A1 => n_188, A2 => n_327, B1 => n_188, B2 => framebuffer_buf_50_3588, ZN => n_176);
  g17509 : MOAI22D0BWP7T port map(A1 => n_188, A2 => n_325, B1 => n_188, B2 => framebuffer_buf_51_3589, ZN => n_175);
  g17510 : MOAI22D0BWP7T port map(A1 => n_188, A2 => n_323, B1 => n_188, B2 => framebuffer_buf_52_3590, ZN => n_174);
  g17511 : MOAI22D0BWP7T port map(A1 => n_188, A2 => n_321, B1 => n_188, B2 => framebuffer_buf_53_3591, ZN => n_173);
  g17512 : MOAI22D0BWP7T port map(A1 => n_171, A2 => n_338, B1 => n_171, B2 => framebuffer_buf_70_3608, ZN => n_172);
  g17513 : MOAI22D0BWP7T port map(A1 => n_171, A2 => n_341, B1 => n_171, B2 => framebuffer_buf_71_3609, ZN => n_170);
  g17514 : MOAI22D0BWP7T port map(A1 => n_249, A2 => n_338, B1 => n_249, B2 => framebuffer_buf_38_3576, ZN => n_169);
  g17515 : MOAI22D0BWP7T port map(A1 => n_249, A2 => n_341, B1 => n_249, B2 => framebuffer_buf_39_3577, ZN => n_168);
  g17516 : MOAI22D0BWP7T port map(A1 => n_171, A2 => n_318, B1 => n_171, B2 => framebuffer_buf_64_3602, ZN => n_167);
  g17517 : MOAI22D0BWP7T port map(A1 => n_171, A2 => n_329, B1 => n_171, B2 => framebuffer_buf_65_3603, ZN => n_166);
  g17518 : MOAI22D0BWP7T port map(A1 => n_171, A2 => n_327, B1 => n_171, B2 => framebuffer_buf_66_3604, ZN => n_165);
  g17519 : MOAI22D0BWP7T port map(A1 => n_171, A2 => n_325, B1 => n_171, B2 => framebuffer_buf_67_3605, ZN => n_164);
  g17520 : MOAI22D0BWP7T port map(A1 => n_171, A2 => n_323, B1 => n_171, B2 => framebuffer_buf_68_3606, ZN => n_163);
  g17521 : MOAI22D0BWP7T port map(A1 => n_171, A2 => n_321, B1 => n_171, B2 => framebuffer_buf_69_3607, ZN => n_162);
  g17522 : MOAI22D0BWP7T port map(A1 => n_249, A2 => n_318, B1 => n_249, B2 => framebuffer_buf_32_3570, ZN => n_161);
  g17523 : MOAI22D0BWP7T port map(A1 => n_249, A2 => n_329, B1 => n_249, B2 => framebuffer_buf_33_3571, ZN => n_160);
  g17524 : MOAI22D0BWP7T port map(A1 => n_249, A2 => n_327, B1 => n_249, B2 => framebuffer_buf_34_3572, ZN => n_159);
  g17559 : MOAI22D0BWP7T port map(A1 => n_180, A2 => n_341, B1 => n_180, B2 => framebuffer_buf_31_3569, ZN => n_158);
  new_framebuffer_buf_reg_153 : LHQD1BWP7T port map(E => n_301, D => n_110, Q => new_framebuffer_buf(153));
  new_framebuffer_buf_reg_154 : LHQD1BWP7T port map(E => n_301, D => n_111, Q => new_framebuffer_buf(154));
  new_framebuffer_buf_reg_155 : LHQD1BWP7T port map(E => n_301, D => n_108, Q => new_framebuffer_buf(155));
  new_framebuffer_buf_reg_156 : LHQD1BWP7T port map(E => n_301, D => n_113, Q => new_framebuffer_buf(156));
  new_framebuffer_buf_reg_157 : LHQD1BWP7T port map(E => n_301, D => n_107, Q => new_framebuffer_buf(157));
  g17537 : OAI21D0BWP7T port map(A1 => n_156, A2 => counter(2), B => n_155, ZN => n_157);
  new_framebuffer_buf_reg_142 : LHQD1BWP7T port map(E => n_301, D => n_101, Q => new_framebuffer_buf(142));
  g17597 : MOAI22D0BWP7T port map(A1 => n_273, A2 => n_341, B1 => n_273, B2 => framebuffer_buf_127_3665, ZN => n_154);
  new_framebuffer_buf_reg_143 : LHQD1BWP7T port map(E => n_301, D => n_103, Q => new_framebuffer_buf(143));
  new_framebuffer_buf_reg_150 : LHQD1BWP7T port map(E => n_301, D => n_120, Q => new_framebuffer_buf(150));
  new_framebuffer_buf_reg_151 : LHQD1BWP7T port map(E => n_301, D => n_89, Q => new_framebuffer_buf(151));
  new_framebuffer_buf_reg_136 : LHQD1BWP7T port map(E => n_301, D => n_87, Q => new_framebuffer_buf(136));
  new_framebuffer_buf_reg_137 : LHQD1BWP7T port map(E => n_301, D => n_85, Q => new_framebuffer_buf(137));
  new_framebuffer_buf_reg_139 : LHQD1BWP7T port map(E => n_301, D => n_79, Q => new_framebuffer_buf(139));
  new_framebuffer_buf_reg_138 : LHQD1BWP7T port map(E => n_301, D => n_84, Q => new_framebuffer_buf(138));
  new_framebuffer_buf_reg_140 : LHQD1BWP7T port map(E => n_301, D => n_83, Q => new_framebuffer_buf(140));
  g17502 : MOAI22D0BWP7T port map(A1 => n_221, A2 => n_327, B1 => n_221, B2 => framebuffer_buf_42_3580, ZN => n_153);
  new_framebuffer_buf_reg_144 : LHQD1BWP7T port map(E => n_301, D => n_81, Q => new_framebuffer_buf(144));
  new_framebuffer_buf_reg_145 : LHQD1BWP7T port map(E => n_301, D => n_90, Q => new_framebuffer_buf(145));
  new_framebuffer_buf_reg_146 : LHQD1BWP7T port map(E => n_301, D => n_91, Q => new_framebuffer_buf(146));
  g17566 : MOAI22D0BWP7T port map(A1 => n_180, A2 => n_318, B1 => n_180, B2 => framebuffer_buf_24_3562, ZN => n_152);
  new_framebuffer_buf_reg_147 : LHQD1BWP7T port map(E => n_301, D => n_80, Q => new_framebuffer_buf(147));
  new_framebuffer_buf_reg_148 : LHQD1BWP7T port map(E => n_301, D => n_100, Q => new_framebuffer_buf(148));
  g17567 : MOAI22D0BWP7T port map(A1 => n_180, A2 => n_329, B1 => n_180, B2 => framebuffer_buf_25_3563, ZN => n_151);
  new_framebuffer_buf_reg_149 : LHQD1BWP7T port map(E => n_301, D => n_99, Q => new_framebuffer_buf(149));
  g17568 : MOAI22D0BWP7T port map(A1 => n_180, A2 => n_327, B1 => n_180, B2 => framebuffer_buf_26_3564, ZN => n_150);
  new_framebuffer_buf_reg_134 : LHQD1BWP7T port map(E => n_301, D => n_98, Q => new_framebuffer_buf(134));
  g17569 : MOAI22D0BWP7T port map(A1 => n_180, A2 => n_325, B1 => n_180, B2 => framebuffer_buf_27_3565, ZN => n_149);
  new_framebuffer_buf_reg_135 : LHQD1BWP7T port map(E => n_301, D => n_96, Q => new_framebuffer_buf(135));
  g17570 : MOAI22D0BWP7T port map(A1 => n_180, A2 => n_323, B1 => n_180, B2 => framebuffer_buf_28_3566, ZN => n_148);
  new_framebuffer_buf_reg_128 : LHQD1BWP7T port map(E => n_301, D => n_76, Q => new_framebuffer_buf(128));
  new_framebuffer_buf_reg_130 : LHQD1BWP7T port map(E => n_301, D => n_78, Q => new_framebuffer_buf(130));
  g17571 : MOAI22D0BWP7T port map(A1 => n_180, A2 => n_321, B1 => n_180, B2 => framebuffer_buf_29_3567, ZN => n_147);
  new_framebuffer_buf_reg_131 : LHQD1BWP7T port map(E => n_301, D => n_88, Q => new_framebuffer_buf(131));
  new_framebuffer_buf_reg_132 : LHQD1BWP7T port map(E => n_301, D => n_86, Q => new_framebuffer_buf(132));
  new_framebuffer_buf_reg_129 : LHQD1BWP7T port map(E => n_301, D => n_77, Q => new_framebuffer_buf(129));
  new_framebuffer_buf_reg_133 : LHQD1BWP7T port map(E => n_301, D => n_92, Q => new_framebuffer_buf(133));
  g17574 : MOAI22D0BWP7T port map(A1 => n_145, A2 => n_338, B1 => n_145, B2 => framebuffer_buf_22_3560, ZN => n_146);
  g17575 : MOAI22D0BWP7T port map(A1 => n_145, A2 => n_341, B1 => n_145, B2 => framebuffer_buf_23_3561, ZN => n_144);
  g17596 : MOAI22D0BWP7T port map(A1 => n_273, A2 => n_338, B1 => n_273, B2 => framebuffer_buf_126_3664, ZN => n_143);
  g17579 : MOAI22D0BWP7T port map(A1 => n_273, A2 => n_323, B1 => n_273, B2 => framebuffer_buf_124_3662, ZN => n_142);
  g17582 : MOAI22D0BWP7T port map(A1 => n_145, A2 => n_318, B1 => n_145, B2 => framebuffer_buf_16_3554, ZN => n_141);
  g17583 : MOAI22D0BWP7T port map(A1 => n_145, A2 => n_329, B1 => n_145, B2 => framebuffer_buf_17_3555, ZN => n_140);
  g17584 : MOAI22D0BWP7T port map(A1 => n_145, A2 => n_327, B1 => n_145, B2 => framebuffer_buf_18_3556, ZN => n_139);
  g17585 : MOAI22D0BWP7T port map(A1 => n_145, A2 => n_325, B1 => n_145, B2 => framebuffer_buf_19_3557, ZN => n_138);
  g17586 : MOAI22D0BWP7T port map(A1 => n_145, A2 => n_323, B1 => n_145, B2 => framebuffer_buf_20_3558, ZN => n_137);
  g17587 : MOAI22D0BWP7T port map(A1 => n_145, A2 => n_321, B1 => n_145, B2 => framebuffer_buf_21_3559, ZN => n_136);
  g17588 : MOAI22D0BWP7T port map(A1 => n_134, A2 => n_338, B1 => n_134, B2 => framebuffer_buf_6_3544, ZN => n_135);
  g17589 : MOAI22D0BWP7T port map(A1 => n_134, A2 => n_341, B1 => n_134, B2 => framebuffer_buf_7_3545, ZN => n_133);
  g17590 : MOAI22D0BWP7T port map(A1 => n_134, A2 => n_318, B1 => n_134, B2 => framebuffer_buf_0_3538, ZN => n_132);
  g17591 : MOAI22D0BWP7T port map(A1 => n_134, A2 => n_329, B1 => n_134, B2 => framebuffer_buf_1_3539, ZN => n_131);
  g17592 : MOAI22D0BWP7T port map(A1 => n_134, A2 => n_327, B1 => n_134, B2 => framebuffer_buf_2_3540, ZN => n_130);
  g17593 : MOAI22D0BWP7T port map(A1 => n_134, A2 => n_325, B1 => n_134, B2 => framebuffer_buf_3_3541, ZN => n_129);
  g17594 : MOAI22D0BWP7T port map(A1 => n_134, A2 => n_323, B1 => n_134, B2 => framebuffer_buf_4_3542, ZN => n_128);
  g17595 : MOAI22D0BWP7T port map(A1 => n_134, A2 => n_321, B1 => n_134, B2 => framebuffer_buf_5_3543, ZN => n_127);
  g17576 : OAI21D0BWP7T port map(A1 => n_156, A2 => counter(4), B => n_126, ZN => n_298);
  g17361 : IND4D0BWP7T port map(A1 => n_1484, B1 => n_276, B2 => n_297, B3 => n_62, ZN => n_351);
  g17461 : NR4D0BWP7T port map(A1 => n_105, A2 => n_57, A3 => n_18, A4 => n_117, ZN => n_125);
  sqi_data_out_reg_6 : LHD1BWP7T port map(E => n_124, D => n_44, Q => UNCONNECTED, QN => n_369);
  sqi_data_out_reg_7 : LHD1BWP7T port map(E => n_124, D => n_30, Q => UNCONNECTED0, QN => n_368);
  sqi_data_out_reg_0 : LHD1BWP7T port map(E => n_124, D => n_24, Q => UNCONNECTED1, QN => n_367);
  sqi_data_out_reg_5 : LHD1BWP7T port map(E => n_124, D => n_45, Q => UNCONNECTED2, QN => n_366);
  sqi_data_out_reg_1 : LHD1BWP7T port map(E => n_124, D => n_39, Q => UNCONNECTED3, QN => n_365);
  g17598 : AOI22D0BWP7T port map(A1 => n_114, A2 => counter(1), B1 => n_122, B2 => n_71, ZN => n_123);
  sqi_data_out_reg_3 : LHD1BWP7T port map(E => n_124, D => n_40, Q => UNCONNECTED4, QN => n_363);
  sqi_data_out_reg_2 : LHD1BWP7T port map(E => n_124, D => n_38, Q => UNCONNECTED5, QN => n_362);
  sqi_data_out_reg_4 : LHD1BWP7T port map(E => n_124, D => n_41, Q => UNCONNECTED6, QN => n_364);
  g17686 : INVD0BWP7T port map(I => n_1483, ZN => n_285);
  g17577 : INR2D0BWP7T port map(A1 => n_292, B1 => n_1484, ZN => n_286);
  state_reg_2 : DFQD1BWP7T port map(CP => clk, D => n_64, Q => state(2));
  g17542 : MOAI22D0BWP7T port map(A1 => n_119, A2 => n_338, B1 => n_119, B2 => framebuffer_buf_150_3688, ZN => n_120);
  g17455 : NR4D0BWP7T port map(A1 => n_54, A2 => n_29, A3 => n_63, A4 => n_117, ZN => n_118);
  g17629 : INVD0BWP7T port map(I => n_1484, ZN => n_116);
  g17632 : ND2D0BWP7T port map(A1 => n_114, A2 => counter(0), ZN => n_115);
  g17657 : MOAI22D0BWP7T port map(A1 => n_112, A2 => n_323, B1 => n_112, B2 => framebuffer_buf_156_3694, ZN => n_113);
  g17658 : MOAI22D0BWP7T port map(A1 => n_112, A2 => n_327, B1 => n_112, B2 => framebuffer_buf_154_3692, ZN => n_111);
  g17659 : MOAI22D0BWP7T port map(A1 => n_112, A2 => n_329, B1 => n_112, B2 => framebuffer_buf_153_3691, ZN => n_110);
  g17660 : MOAI22D0BWP7T port map(A1 => n_112, A2 => n_318, B1 => n_112, B2 => framebuffer_buf_152_3690, ZN => n_109);
  g17661 : MOAI22D0BWP7T port map(A1 => n_112, A2 => n_325, B1 => n_112, B2 => framebuffer_buf_155_3693, ZN => n_108);
  g17662 : MOAI22D0BWP7T port map(A1 => n_112, A2 => n_321, B1 => n_112, B2 => framebuffer_buf_157_3695, ZN => n_107);
  g17453 : NR3D0BWP7T port map(A1 => n_105, A2 => n_52, A3 => n_104, ZN => n_106);
  g17541 : MOAI22D0BWP7T port map(A1 => n_102, A2 => n_341, B1 => n_102, B2 => framebuffer_buf_143_3681, ZN => n_103);
  g17540 : MOAI22D0BWP7T port map(A1 => n_102, A2 => n_338, B1 => n_102, B2 => framebuffer_buf_142_3680, ZN => n_101);
  g17529 : MOAI22D0BWP7T port map(A1 => n_119, A2 => n_323, B1 => n_119, B2 => framebuffer_buf_148_3686, ZN => n_100);
  g17555 : MOAI22D0BWP7T port map(A1 => n_119, A2 => n_321, B1 => n_119, B2 => framebuffer_buf_149_3687, ZN => n_99);
  g17556 : MOAI22D0BWP7T port map(A1 => n_97, A2 => n_338, B1 => n_97, B2 => framebuffer_buf_134_3672, ZN => n_98);
  g17557 : MOAI22D0BWP7T port map(A1 => n_97, A2 => n_341, B1 => n_97, B2 => framebuffer_buf_135_3673, ZN => n_96);
  g17664 : AOI21D0BWP7T port map(A1 => n_122, A2 => n_95, B => n_114, ZN => n_155);
  g17688 : INVD0BWP7T port map(I => n_145, ZN => n_184);
  g17687 : INVD0BWP7T port map(I => n_134, ZN => n_186);
  g17663 : IAO21D0BWP7T port map(A1 => n_156, A2 => n_56, B => n_114, ZN => n_126);
  g17679 : IND2D0BWP7T port map(A1 => n_94, B1 => counter(4), ZN => n_305);
  g17565 : MOAI22D0BWP7T port map(A1 => n_97, A2 => n_321, B1 => n_97, B2 => framebuffer_buf_133_3671, ZN => n_92);
  g17544 : MOAI22D0BWP7T port map(A1 => n_119, A2 => n_327, B1 => n_119, B2 => framebuffer_buf_146_3684, ZN => n_91);
  g17545 : MOAI22D0BWP7T port map(A1 => n_119, A2 => n_329, B1 => n_119, B2 => framebuffer_buf_145_3683, ZN => n_90);
  g17543 : MOAI22D0BWP7T port map(A1 => n_119, A2 => n_341, B1 => n_119, B2 => framebuffer_buf_151_3689, ZN => n_89);
  g17564 : MOAI22D0BWP7T port map(A1 => n_97, A2 => n_325, B1 => n_97, B2 => framebuffer_buf_131_3669, ZN => n_88);
  g17547 : MOAI22D0BWP7T port map(A1 => n_102, A2 => n_318, B1 => n_102, B2 => framebuffer_buf_136_3674, ZN => n_87);
  g17560 : MOAI22D0BWP7T port map(A1 => n_97, A2 => n_323, B1 => n_97, B2 => framebuffer_buf_132_3670, ZN => n_86);
  g17548 : MOAI22D0BWP7T port map(A1 => n_102, A2 => n_329, B1 => n_102, B2 => framebuffer_buf_137_3675, ZN => n_85);
  g17549 : MOAI22D0BWP7T port map(A1 => n_102, A2 => n_327, B1 => n_102, B2 => framebuffer_buf_138_3676, ZN => n_84);
  g17550 : MOAI22D0BWP7T port map(A1 => n_102, A2 => n_323, B1 => n_102, B2 => framebuffer_buf_140_3678, ZN => n_83);
  g17551 : MOAI22D0BWP7T port map(A1 => n_102, A2 => n_321, B1 => n_102, B2 => framebuffer_buf_141_3679, ZN => n_82);
  g17552 : MOAI22D0BWP7T port map(A1 => n_119, A2 => n_318, B1 => n_119, B2 => framebuffer_buf_144_3682, ZN => n_81);
  g17553 : MOAI22D0BWP7T port map(A1 => n_119, A2 => n_325, B1 => n_119, B2 => framebuffer_buf_147_3685, ZN => n_80);
  g17546 : MOAI22D0BWP7T port map(A1 => n_102, A2 => n_325, B1 => n_102, B2 => framebuffer_buf_139_3677, ZN => n_79);
  g17563 : MOAI22D0BWP7T port map(A1 => n_97, A2 => n_327, B1 => n_97, B2 => framebuffer_buf_130_3668, ZN => n_78);
  g17562 : MOAI22D0BWP7T port map(A1 => n_97, A2 => n_329, B1 => n_97, B2 => framebuffer_buf_129_3667, ZN => n_77);
  g17561 : MOAI22D0BWP7T port map(A1 => n_97, A2 => n_318, B1 => n_97, B2 => framebuffer_buf_128_3666, ZN => n_76);
  row_buf_reg_5 : DFXQD1BWP7T port map(CP => clk, DA => new_row_buf(5), DB => row_buf(5), SA => n_355, Q => row_buf(5));
  row_buf_reg_0 : DFXQD1BWP7T port map(CP => clk, DA => new_row_buf(0), DB => row_buf(0), SA => n_355, Q => row_buf(0));
  row_buf_reg_2 : DFXQD1BWP7T port map(CP => clk, DA => new_row_buf(2), DB => row_buf(2), SA => n_355, Q => row_buf(2));
  row_buf_reg_4 : DFXQD1BWP7T port map(CP => clk, DA => new_row_buf(4), DB => row_buf(4), SA => n_355, Q => row_buf(4));
  row_buf_reg_3 : DFXQD1BWP7T port map(CP => clk, DA => new_row_buf(3), DB => row_buf(3), SA => n_355, Q => row_buf(3));
  row_buf_reg_1 : DFXQD1BWP7T port map(CP => clk, DA => new_row_buf(1), DB => row_buf(1), SA => n_355, Q => row_buf(1));
  g17656 : NR4D0BWP7T port map(A1 => n_290, A2 => n_95, A3 => n_74, A4 => counter(3), ZN => n_75);
  g17672 : ND2D0BWP7T port map(A1 => n_70, A2 => n_71, ZN => n_211);
  g17669 : IND2D0BWP7T port map(A1 => n_93, B1 => n_69, ZN => n_221);
  g17670 : ND2D0BWP7T port map(A1 => n_70, A2 => n_68, ZN => n_229);
  g17671 : IND2D0BWP7T port map(A1 => n_93, B1 => n_70, ZN => n_214);
  g17655 : ND2D0BWP7T port map(A1 => n_70, A2 => n_67, ZN => n_171);
  g17673 : ND2D0BWP7T port map(A1 => n_69, A2 => n_71, ZN => n_188);
  g17674 : ND2D0BWP7T port map(A1 => n_69, A2 => n_68, ZN => n_217);
  g17654 : ND2D0BWP7T port map(A1 => n_69, A2 => n_67, ZN => n_249);
  g17675 : INVD0BWP7T port map(I => n_65, ZN => n_66);
  g17536 : ND4D0BWP7T port map(A1 => n_61, A2 => n_389, A3 => n_55, A4 => n_355, ZN => n_64);
  g17693 : IND2D0BWP7T port map(A1 => n_63, B1 => n_73, ZN => n_124);
  g17578 : ND3D0BWP7T port map(A1 => n_62, A2 => n_61, A3 => n_156, ZN => n_354);
  g17694 : ND2D0BWP7T port map(A1 => n_59, A2 => n_68, ZN => n_180);
  g17681 : ND2D0BWP7T port map(A1 => n_60, A2 => n_71, ZN => n_262);
  g17695 : ND2D0BWP7T port map(A1 => n_60, A2 => n_68, ZN => n_273);
  g17682 : IND2D0BWP7T port map(A1 => n_93, B1 => n_60, ZN => n_268);
  g17685 : ND2D0BWP7T port map(A1 => n_60, A2 => n_67, ZN => n_266);
  g17698 : ND2D0BWP7T port map(A1 => n_59, A2 => n_71, ZN => n_145);
  g17697 : ND2D0BWP7T port map(A1 => n_59, A2 => n_67, ZN => n_134);
  g17678 : NR2D0BWP7T port map(A1 => n_35, A2 => counter(4), ZN => n_65);
  g17665 : OAI22D0BWP7T port map(A1 => n_53, A2 => n_292, B1 => n_49, B2 => n_16, ZN => n_105);
  g17689 : OAI211D1BWP7T port map(A1 => sqi_finished, A2 => n_32, B => n_50, C => n_26, ZN => n_57);
  g17704 : IND2D0BWP7T port map(A1 => n_290, B1 => n_56, ZN => n_94);
  g17691 : OAI211D0BWP7T port map(A1 => sqi_finished, A2 => n_156, B => n_72, C => n_292, ZN => n_114);
  g17699 : AOI21D0BWP7T port map(A1 => n_36, A2 => n_37, B => n_55, ZN => n_301);
  g17676 : NR2D0BWP7T port map(A1 => n_53, A2 => n_292, ZN => n_54);
  g17702 : OAI21D0BWP7T port map(A1 => n_51, A2 => n_25, B => n_50, ZN => n_52);
  g17705 : OAI21D0BWP7T port map(A1 => n_49, A2 => n_17, B => n_48, ZN => n_63);
  g17677 : IND2D0BWP7T port map(A1 => n_292, B1 => n_53, ZN => n_62);
  g17692 : NR3D0BWP7T port map(A1 => n_47, A2 => n_74, A3 => counter(3), ZN => n_69);
  g17690 : NR3D0BWP7T port map(A1 => n_47, A2 => n_1, A3 => counter(2), ZN => n_70);
  g17684 : IND2D0BWP7T port map(A1 => n_46, B1 => n_67, ZN => n_97);
  g17683 : IND2D0BWP7T port map(A1 => n_46, B1 => n_71, ZN => n_119);
  g17680 : OR2D0BWP7T port map(A1 => n_46, A2 => n_93, Z => n_102);
  g17714 : AO22D0BWP7T port map(A1 => n_43, A2 => calc_buf_in(4), B1 => row_buf(5), B2 => n_42, Z => n_45);
  g17713 : AO22D0BWP7T port map(A1 => n_43, A2 => calc_buf_in(5), B1 => calc_buf_in(0), B2 => n_42, Z => n_44);
  g17709 : AO22D0BWP7T port map(A1 => n_43, A2 => calc_buf_in(3), B1 => row_buf(4), B2 => n_42, Z => n_41);
  g17710 : AO22D0BWP7T port map(A1 => n_43, A2 => calc_buf_in(2), B1 => row_buf(3), B2 => n_42, Z => n_40);
  g17711 : AO22D0BWP7T port map(A1 => n_43, A2 => calc_buf_in(0), B1 => row_buf(1), B2 => n_42, Z => n_39);
  g17712 : AO22D0BWP7T port map(A1 => n_43, A2 => calc_buf_in(1), B1 => row_buf(2), B2 => n_42, Z => n_38);
  g17707 : NR2D0BWP7T port map(A1 => n_47, A2 => n_8, ZN => n_60);
  g17708 : INR2D0BWP7T port map(A1 => n_14, B1 => n_47, ZN => n_59);
  g17716 : OAI21D0BWP7T port map(A1 => n_37, A2 => n_68, B => n_36, ZN => n_112);
  new_row_buf_reg_0 : LHQD1BWP7T port map(E => n_34, D => sqi_data_in(0), Q => new_row_buf(0));
  g17701 : IND4D0BWP7T port map(A1 => n_37, B1 => n_4, B2 => n_3, B3 => n_67, ZN => n_35);
  new_row_buf_reg_1 : LHQD1BWP7T port map(E => n_34, D => sqi_data_in(1), Q => new_row_buf(1));
  g17723 : AN2D1BWP7T port map(A1 => n_32, A2 => n_51, Z => n_33);
  g17715 : MAOI22D0BWP7T port map(A1 => n_11, A2 => ce, B1 => n_72, B2 => n_23, ZN => n_61);
  new_row_buf_reg_5 : LHQD1BWP7T port map(E => n_34, D => sqi_data_in(5), Q => new_row_buf(5));
  new_row_buf_reg_3 : LHQD1BWP7T port map(E => n_34, D => sqi_data_in(3), Q => new_row_buf(3));
  new_row_buf_reg_2 : LHQD1BWP7T port map(E => n_34, D => sqi_data_in(2), Q => new_row_buf(2));
  new_row_buf_reg_4 : LHQD1BWP7T port map(E => n_34, D => sqi_data_in(4), Q => new_row_buf(4));
  g17733 : ND2D0BWP7T port map(A1 => n_122, A2 => sqi_finished, ZN => n_290);
  g17727 : INR2D0BWP7T port map(A1 => calc_buf_in(1), B1 => n_73, ZN => n_30);
  g17726 : OAI22D0BWP7T port map(A1 => n_55, A2 => sqi_finished, B1 => n_28, B2 => rw, ZN => n_29);
  g17728 : AO21D0BWP7T port map(A1 => n_19, A2 => n_297, B => n_25, Z => n_26);
  g17706 : IND3D0BWP7T port map(A1 => n_37, B1 => sqi_finished, B2 => counter(4), ZN => n_46);
  g17703 : NR3D0BWP7T port map(A1 => n_37, A2 => n_68, A3 => counter(4), ZN => n_53);
  g17724 : INR2D0BWP7T port map(A1 => row_buf(0), B1 => n_73, ZN => n_24);
  g17730 : NR2D0BWP7T port map(A1 => n_22, A2 => n_25, ZN => n_36);
  g17731 : IND2D1BWP7T port map(A1 => n_72, B1 => n_23, ZN => n_50);
  g17729 : OAI22D0BWP7T port map(A1 => n_21, A2 => n_25, B1 => n_28, B2 => ce, ZN => n_104);
  g17732 : ND2D0BWP7T port map(A1 => n_22, A2 => sqi_finished, ZN => n_47);
  g17735 : INVD0BWP7T port map(I => n_122, ZN => n_156);
  g17736 : CKAN2D1BWP7T port map(A1 => n_21, A2 => n_20, Z => n_32);
  g17737 : INR2D0BWP7T port map(A1 => n_19, B1 => n_18, ZN => n_51);
  g17739 : NR2D0BWP7T port map(A1 => n_20, A2 => n_25, ZN => n_34);
  g17740 : ND2D0BWP7T port map(A1 => n_49, A2 => n_48, ZN => n_43);
  g17742 : CKND0BWP7T port map(I => n_16, ZN => n_17);
  g17744 : ND2D4BWP7T port map(A1 => n_28, A2 => n_276, ZN => ready);
  g17741 : ND2D0BWP7T port map(A1 => n_297, A2 => n_55, ZN => n_122);
  g17743 : INVD0BWP7T port map(I => n_73, ZN => n_42);
  g17746 : NR4D0BWP7T port map(A1 => n_2, A2 => x(4), A3 => x(0), A4 => x(1), ZN => n_16);
  g17745 : INR2D0BWP7T port map(A1 => n_12, B1 => counter(4), ZN => n_22);
  g17747 : OAI21D0BWP7T port map(A1 => n_14, A2 => n_13, B => n_12, ZN => n_23);
  g17751 : INVD0BWP7T port map(I => n_297, ZN => n_185);
  g17750 : INVD0BWP7T port map(I => n_28, ZN => n_11);
  g17748 : IND3D1BWP7T port map(A1 => state(3), B1 => state(2), B2 => n_10, ZN => n_72);
  g17738 : ND2D1BWP7T port map(A1 => n_12, A2 => n_14, ZN => n_37);
  g17749 : IND3D1BWP7T port map(A1 => state(2), B1 => state(3), B2 => n_10, ZN => n_73);
  g17754 : ND2D1BWP7T port map(A1 => n_6, A2 => n_9, ZN => n_19);
  g17752 : ND2D1BWP7T port map(A1 => n_7, A2 => n_9, ZN => n_21);
  g17753 : NR2D0BWP7T port map(A1 => n_8, A2 => n_95, ZN => n_56);
  g17756 : ND2D1BWP7T port map(A1 => n_7, A2 => state(3), ZN => n_20);
  g17755 : ND2D1BWP7T port map(A1 => n_6, A2 => state(3), ZN => n_48);
  g17757 : IND2D1BWP7T port map(A1 => n_5, B1 => state(3), ZN => n_28);
  g17763 : NR2D1BWP7T port map(A1 => n_276, A2 => reset, ZN => n_117);
  g17762 : INR2D1BWP7T port map(A1 => n_9, B1 => n_5, ZN => n_18);
  g17764 : IND2D1BWP7T port map(A1 => n_5, B1 => state(2), ZN => n_49);
  g17766 : ND2D1BWP7T port map(A1 => n_6, A2 => state(2), ZN => n_55);
  g17758 : ND2D1BWP7T port map(A1 => n_7, A2 => state(2), ZN => n_292);
  g17759 : CKND2D1BWP7T port map(A1 => n_10, A2 => n_9, ZN => n_297);
  g17760 : NR4D0BWP7T port map(A1 => y(5), A2 => y(4), A3 => y(6), A4 => y(7), ZN => n_4);
  g17761 : NR4D0BWP7T port map(A1 => y(1), A2 => y(0), A3 => y(2), A4 => y(3), ZN => n_3);
  g17765 : NR3D0BWP7T port map(A1 => counter(5), A2 => counter(6), A3 => counter(7), ZN => n_12);
  g17773 : INVD1BWP7T port map(I => n_95, ZN => n_68);
  g17774 : OR2D1BWP7T port map(A1 => x(2), A2 => x(3), Z => n_2);
  g17767 : ND2D0BWP7T port map(A1 => counter(3), A2 => counter(2), ZN => n_8);
  g17777 : ND2D1BWP7T port map(A1 => state(1), A2 => state(0), ZN => n_5);
  g17770 : NR2D1BWP7T port map(A1 => state(2), A2 => state(3), ZN => n_9);
  g17780 : CKND2D1BWP7T port map(A1 => counter(0), A2 => counter(1), ZN => n_95);
  g17769 : NR2D1BWP7T port map(A1 => state(1), A2 => state(0), ZN => n_10);
  g17776 : NR2XD0BWP7T port map(A1 => counter(2), A2 => counter(3), ZN => n_14);
  g17775 : INR2D1BWP7T port map(A1 => state(1), B1 => state(0), ZN => n_7);
  g17768 : INR2D1BWP7T port map(A1 => state(0), B1 => state(1), ZN => n_6);
  g17778 : NR2D0BWP7T port map(A1 => counter(1), A2 => counter(0), ZN => n_67);
  g17771 : ND2D1BWP7T port map(A1 => state(3), A2 => state(2), ZN => n_276);
  g17772 : IND2D0BWP7T port map(A1 => counter(1), B1 => counter(0), ZN => n_93);
  g17779 : INR2D0BWP7T port map(A1 => counter(1), B1 => counter(0), ZN => n_71);
  g17799 : INVD1BWP7T port map(I => reset, ZN => n_347);
  g17802 : INVD1BWP7T port map(I => reset, ZN => n_349);
  g17803 : INVD1BWP7T port map(I => reset, ZN => n_357);
  g17792 : INVD0BWP7T port map(I => sqi_data_in(1), ZN => n_329);
  g17787 : INVD0BWP7T port map(I => sqi_data_in(3), ZN => n_325);
  g17798 : INVD1BWP7T port map(I => reset, ZN => n_355);
  g17794 : INVD1BWP7T port map(I => reset, ZN => n_360);
  g17783 : CKND1BWP7T port map(I => sqi_finished, ZN => n_25);
  g17785 : INVD0BWP7T port map(I => sqi_data_in(7), ZN => n_341);
  g17784 : INVD0BWP7T port map(I => sqi_data_in(6), ZN => n_338);
  g17791 : INVD0BWP7T port map(I => sqi_data_in(2), ZN => n_327);
  g17786 : INVD0BWP7T port map(I => sqi_data_in(4), ZN => n_323);
  g17793 : INVD0BWP7T port map(I => sqi_data_in(5), ZN => n_321);
  g17788 : INVD0BWP7T port map(I => sqi_data_in(0), ZN => n_318);
  g17795 : INVD1BWP7T port map(I => reset, ZN => n_356);
  g2 : ND2D1BWP7T port map(A1 => n_185, A2 => sqi_finished, ZN => n_389);
  drc_bufs18209 : INVD4BWP7T port map(I => n_392, ZN => calc_buf_out(0));
  drc_bufs18215 : INVD4BWP7T port map(I => n_398, ZN => framebuffer_buf(157));
  drc_bufs18221 : INVD4BWP7T port map(I => n_404, ZN => framebuffer_buf(156));
  drc_bufs18227 : INVD4BWP7T port map(I => n_410, ZN => framebuffer_buf(155));
  drc_bufs18233 : INVD4BWP7T port map(I => n_416, ZN => framebuffer_buf(154));
  drc_bufs18239 : INVD4BWP7T port map(I => n_422, ZN => framebuffer_buf(153));
  drc_bufs18245 : INVD4BWP7T port map(I => n_428, ZN => framebuffer_buf(152));
  drc_bufs18251 : INVD4BWP7T port map(I => n_434, ZN => framebuffer_buf(151));
  drc_bufs18257 : INVD4BWP7T port map(I => n_440, ZN => framebuffer_buf(150));
  drc_bufs18263 : INVD4BWP7T port map(I => n_446, ZN => framebuffer_buf(149));
  drc_bufs18269 : INVD4BWP7T port map(I => n_452, ZN => framebuffer_buf(148));
  drc_bufs18275 : INVD4BWP7T port map(I => n_458, ZN => framebuffer_buf(147));
  drc_bufs18281 : INVD4BWP7T port map(I => n_464, ZN => framebuffer_buf(146));
  drc_bufs18287 : INVD4BWP7T port map(I => n_470, ZN => framebuffer_buf(145));
  drc_bufs18293 : INVD4BWP7T port map(I => n_476, ZN => framebuffer_buf(144));
  drc_bufs18299 : INVD4BWP7T port map(I => n_482, ZN => framebuffer_buf(143));
  drc_bufs18305 : INVD4BWP7T port map(I => n_488, ZN => framebuffer_buf(142));
  drc_bufs18311 : INVD4BWP7T port map(I => n_494, ZN => framebuffer_buf(141));
  drc_bufs18317 : INVD4BWP7T port map(I => n_500, ZN => framebuffer_buf(140));
  drc_bufs18323 : INVD4BWP7T port map(I => n_506, ZN => framebuffer_buf(139));
  drc_bufs18329 : INVD4BWP7T port map(I => n_512, ZN => framebuffer_buf(138));
  drc_bufs18335 : INVD4BWP7T port map(I => n_518, ZN => framebuffer_buf(137));
  drc_bufs18341 : INVD4BWP7T port map(I => n_524, ZN => framebuffer_buf(136));
  drc_bufs18347 : INVD4BWP7T port map(I => n_530, ZN => framebuffer_buf(135));
  drc_bufs18353 : INVD4BWP7T port map(I => n_536, ZN => framebuffer_buf(134));
  drc_bufs18359 : INVD4BWP7T port map(I => n_542, ZN => framebuffer_buf(133));
  drc_bufs18365 : INVD4BWP7T port map(I => n_548, ZN => framebuffer_buf(132));
  drc_bufs18371 : INVD4BWP7T port map(I => n_554, ZN => framebuffer_buf(131));
  drc_bufs18377 : INVD4BWP7T port map(I => n_560, ZN => framebuffer_buf(130));
  drc_bufs18383 : INVD4BWP7T port map(I => n_566, ZN => framebuffer_buf(129));
  drc_bufs18389 : INVD4BWP7T port map(I => n_572, ZN => framebuffer_buf(128));
  drc_bufs18395 : INVD4BWP7T port map(I => n_578, ZN => framebuffer_buf(127));
  drc_bufs18401 : INVD4BWP7T port map(I => n_584, ZN => framebuffer_buf(126));
  drc_bufs18407 : INVD4BWP7T port map(I => n_590, ZN => framebuffer_buf(125));
  drc_bufs18413 : INVD4BWP7T port map(I => n_596, ZN => framebuffer_buf(124));
  drc_bufs18419 : INVD4BWP7T port map(I => n_602, ZN => framebuffer_buf(123));
  drc_bufs18425 : INVD4BWP7T port map(I => n_608, ZN => framebuffer_buf(122));
  drc_bufs18431 : INVD4BWP7T port map(I => n_614, ZN => framebuffer_buf(121));
  drc_bufs18437 : INVD4BWP7T port map(I => n_620, ZN => framebuffer_buf(120));
  drc_bufs18443 : INVD4BWP7T port map(I => n_626, ZN => framebuffer_buf(119));
  drc_bufs18449 : INVD4BWP7T port map(I => n_632, ZN => framebuffer_buf(118));
  drc_bufs18455 : INVD4BWP7T port map(I => n_638, ZN => framebuffer_buf(117));
  drc_bufs18461 : INVD4BWP7T port map(I => n_644, ZN => framebuffer_buf(116));
  drc_bufs18467 : INVD4BWP7T port map(I => n_650, ZN => framebuffer_buf(115));
  drc_bufs18473 : INVD4BWP7T port map(I => n_656, ZN => framebuffer_buf(114));
  drc_bufs18479 : INVD4BWP7T port map(I => n_662, ZN => framebuffer_buf(113));
  drc_bufs18485 : INVD4BWP7T port map(I => n_668, ZN => framebuffer_buf(112));
  drc_bufs18491 : INVD4BWP7T port map(I => n_674, ZN => framebuffer_buf(111));
  drc_bufs18497 : INVD4BWP7T port map(I => n_680, ZN => framebuffer_buf(110));
  drc_bufs18503 : INVD4BWP7T port map(I => n_686, ZN => framebuffer_buf(109));
  drc_bufs18509 : INVD4BWP7T port map(I => n_692, ZN => framebuffer_buf(108));
  drc_bufs18515 : INVD4BWP7T port map(I => n_698, ZN => framebuffer_buf(107));
  drc_bufs18521 : INVD4BWP7T port map(I => n_704, ZN => framebuffer_buf(106));
  drc_bufs18527 : INVD4BWP7T port map(I => n_710, ZN => framebuffer_buf(105));
  drc_bufs18533 : INVD4BWP7T port map(I => n_716, ZN => framebuffer_buf(104));
  drc_bufs18539 : INVD4BWP7T port map(I => n_722, ZN => framebuffer_buf(103));
  drc_bufs18545 : INVD4BWP7T port map(I => n_728, ZN => framebuffer_buf(102));
  drc_bufs18551 : INVD4BWP7T port map(I => n_734, ZN => framebuffer_buf(101));
  drc_bufs18557 : INVD4BWP7T port map(I => n_740, ZN => framebuffer_buf(100));
  drc_bufs18563 : INVD4BWP7T port map(I => n_746, ZN => framebuffer_buf(99));
  drc_bufs18569 : INVD4BWP7T port map(I => n_752, ZN => framebuffer_buf(98));
  drc_bufs18575 : INVD4BWP7T port map(I => n_758, ZN => framebuffer_buf(97));
  drc_bufs18581 : INVD4BWP7T port map(I => n_764, ZN => framebuffer_buf(96));
  drc_bufs18587 : INVD4BWP7T port map(I => n_770, ZN => framebuffer_buf(95));
  drc_bufs18593 : INVD4BWP7T port map(I => n_776, ZN => framebuffer_buf(94));
  drc_bufs18599 : INVD4BWP7T port map(I => n_782, ZN => framebuffer_buf(93));
  drc_bufs18605 : INVD4BWP7T port map(I => n_788, ZN => framebuffer_buf(92));
  drc_bufs18611 : INVD4BWP7T port map(I => n_794, ZN => framebuffer_buf(91));
  drc_bufs18617 : INVD4BWP7T port map(I => n_800, ZN => framebuffer_buf(90));
  drc_bufs18623 : INVD4BWP7T port map(I => n_806, ZN => framebuffer_buf(89));
  drc_bufs18629 : INVD4BWP7T port map(I => n_812, ZN => framebuffer_buf(88));
  drc_bufs18635 : INVD4BWP7T port map(I => n_818, ZN => framebuffer_buf(87));
  drc_bufs18641 : INVD4BWP7T port map(I => n_824, ZN => framebuffer_buf(86));
  drc_bufs18647 : INVD4BWP7T port map(I => n_830, ZN => framebuffer_buf(85));
  drc_bufs18653 : INVD4BWP7T port map(I => n_836, ZN => framebuffer_buf(84));
  drc_bufs18659 : INVD4BWP7T port map(I => n_842, ZN => framebuffer_buf(83));
  drc_bufs18665 : INVD4BWP7T port map(I => n_848, ZN => framebuffer_buf(82));
  drc_bufs18671 : INVD4BWP7T port map(I => n_854, ZN => framebuffer_buf(81));
  drc_bufs18677 : INVD4BWP7T port map(I => n_860, ZN => framebuffer_buf(80));
  drc_bufs18683 : INVD4BWP7T port map(I => n_866, ZN => framebuffer_buf(79));
  drc_bufs18689 : INVD4BWP7T port map(I => n_872, ZN => framebuffer_buf(78));
  drc_bufs18695 : INVD4BWP7T port map(I => n_878, ZN => framebuffer_buf(77));
  drc_bufs18701 : INVD4BWP7T port map(I => n_884, ZN => framebuffer_buf(76));
  drc_bufs18707 : INVD4BWP7T port map(I => n_890, ZN => framebuffer_buf(75));
  drc_bufs18713 : INVD4BWP7T port map(I => n_896, ZN => framebuffer_buf(74));
  drc_bufs18719 : INVD4BWP7T port map(I => n_902, ZN => framebuffer_buf(73));
  drc_bufs18725 : INVD4BWP7T port map(I => n_908, ZN => framebuffer_buf(72));
  drc_bufs18731 : INVD4BWP7T port map(I => n_914, ZN => framebuffer_buf(71));
  drc_bufs18737 : INVD4BWP7T port map(I => n_920, ZN => framebuffer_buf(70));
  drc_bufs18743 : INVD4BWP7T port map(I => n_926, ZN => framebuffer_buf(69));
  drc_bufs18749 : INVD4BWP7T port map(I => n_932, ZN => framebuffer_buf(68));
  drc_bufs18755 : INVD4BWP7T port map(I => n_938, ZN => framebuffer_buf(67));
  drc_bufs18761 : INVD4BWP7T port map(I => n_944, ZN => framebuffer_buf(66));
  drc_bufs18767 : INVD4BWP7T port map(I => n_950, ZN => framebuffer_buf(65));
  drc_bufs18773 : INVD4BWP7T port map(I => n_956, ZN => framebuffer_buf(64));
  drc_bufs18779 : INVD4BWP7T port map(I => n_962, ZN => framebuffer_buf(63));
  drc_bufs18785 : INVD4BWP7T port map(I => n_968, ZN => framebuffer_buf(62));
  drc_bufs18791 : INVD4BWP7T port map(I => n_974, ZN => framebuffer_buf(61));
  drc_bufs18797 : INVD4BWP7T port map(I => n_980, ZN => framebuffer_buf(60));
  drc_bufs18803 : INVD4BWP7T port map(I => n_986, ZN => framebuffer_buf(59));
  drc_bufs18809 : INVD4BWP7T port map(I => n_992, ZN => framebuffer_buf(58));
  drc_bufs18815 : INVD4BWP7T port map(I => n_998, ZN => framebuffer_buf(57));
  drc_bufs18821 : INVD4BWP7T port map(I => n_1004, ZN => framebuffer_buf(56));
  drc_bufs18827 : INVD4BWP7T port map(I => n_1010, ZN => framebuffer_buf(55));
  drc_bufs18833 : INVD4BWP7T port map(I => n_1016, ZN => framebuffer_buf(54));
  drc_bufs18839 : INVD4BWP7T port map(I => n_1022, ZN => framebuffer_buf(53));
  drc_bufs18845 : INVD4BWP7T port map(I => n_1028, ZN => framebuffer_buf(52));
  drc_bufs18851 : INVD4BWP7T port map(I => n_1034, ZN => framebuffer_buf(51));
  drc_bufs18857 : INVD4BWP7T port map(I => n_1040, ZN => framebuffer_buf(50));
  drc_bufs18863 : INVD4BWP7T port map(I => n_1046, ZN => framebuffer_buf(49));
  drc_bufs18869 : INVD4BWP7T port map(I => n_1052, ZN => framebuffer_buf(48));
  drc_bufs18875 : INVD4BWP7T port map(I => n_1058, ZN => framebuffer_buf(47));
  drc_bufs18881 : INVD4BWP7T port map(I => n_1064, ZN => framebuffer_buf(46));
  drc_bufs18887 : INVD4BWP7T port map(I => n_1070, ZN => framebuffer_buf(45));
  drc_bufs18893 : INVD4BWP7T port map(I => n_1076, ZN => framebuffer_buf(44));
  drc_bufs18899 : INVD4BWP7T port map(I => n_1082, ZN => framebuffer_buf(43));
  drc_bufs18905 : INVD4BWP7T port map(I => n_1088, ZN => framebuffer_buf(42));
  drc_bufs18911 : INVD4BWP7T port map(I => n_1094, ZN => framebuffer_buf(41));
  drc_bufs18917 : INVD4BWP7T port map(I => n_1100, ZN => framebuffer_buf(40));
  drc_bufs18923 : INVD4BWP7T port map(I => n_1106, ZN => framebuffer_buf(39));
  drc_bufs18929 : INVD4BWP7T port map(I => n_1112, ZN => framebuffer_buf(38));
  drc_bufs18935 : INVD4BWP7T port map(I => n_1118, ZN => framebuffer_buf(37));
  drc_bufs18941 : INVD4BWP7T port map(I => n_1124, ZN => framebuffer_buf(36));
  drc_bufs18947 : INVD4BWP7T port map(I => n_1130, ZN => framebuffer_buf(35));
  drc_bufs18953 : INVD4BWP7T port map(I => n_1136, ZN => framebuffer_buf(34));
  drc_bufs18959 : INVD4BWP7T port map(I => n_1142, ZN => framebuffer_buf(33));
  drc_bufs18965 : INVD4BWP7T port map(I => n_1148, ZN => framebuffer_buf(32));
  drc_bufs18971 : INVD4BWP7T port map(I => n_1154, ZN => framebuffer_buf(31));
  drc_bufs18977 : INVD4BWP7T port map(I => n_1160, ZN => framebuffer_buf(30));
  drc_bufs18983 : INVD4BWP7T port map(I => n_1166, ZN => framebuffer_buf(29));
  drc_bufs18989 : INVD4BWP7T port map(I => n_1172, ZN => framebuffer_buf(28));
  drc_bufs18995 : INVD4BWP7T port map(I => n_1178, ZN => framebuffer_buf(27));
  drc_bufs19001 : INVD4BWP7T port map(I => n_1184, ZN => framebuffer_buf(26));
  drc_bufs19007 : INVD4BWP7T port map(I => n_1190, ZN => framebuffer_buf(25));
  drc_bufs19013 : INVD4BWP7T port map(I => n_1196, ZN => framebuffer_buf(24));
  drc_bufs19019 : INVD4BWP7T port map(I => n_1202, ZN => framebuffer_buf(23));
  drc_bufs19025 : INVD4BWP7T port map(I => n_1208, ZN => framebuffer_buf(22));
  drc_bufs19031 : INVD4BWP7T port map(I => n_1214, ZN => framebuffer_buf(21));
  drc_bufs19037 : INVD4BWP7T port map(I => n_1220, ZN => framebuffer_buf(20));
  drc_bufs19043 : INVD4BWP7T port map(I => n_1226, ZN => framebuffer_buf(19));
  drc_bufs19049 : INVD4BWP7T port map(I => n_1232, ZN => framebuffer_buf(18));
  drc_bufs19055 : INVD4BWP7T port map(I => n_1238, ZN => framebuffer_buf(17));
  drc_bufs19061 : INVD4BWP7T port map(I => n_1244, ZN => framebuffer_buf(16));
  drc_bufs19067 : INVD4BWP7T port map(I => n_1250, ZN => framebuffer_buf(15));
  drc_bufs19073 : INVD4BWP7T port map(I => n_1256, ZN => framebuffer_buf(14));
  drc_bufs19079 : INVD4BWP7T port map(I => n_1262, ZN => framebuffer_buf(13));
  drc_bufs19085 : INVD4BWP7T port map(I => n_1268, ZN => framebuffer_buf(12));
  drc_bufs19091 : INVD4BWP7T port map(I => n_1274, ZN => framebuffer_buf(11));
  drc_bufs19097 : INVD4BWP7T port map(I => n_1280, ZN => framebuffer_buf(10));
  drc_bufs19103 : INVD4BWP7T port map(I => n_1286, ZN => framebuffer_buf(9));
  drc_bufs19109 : INVD4BWP7T port map(I => n_1292, ZN => framebuffer_buf(8));
  drc_bufs19115 : INVD4BWP7T port map(I => n_1298, ZN => framebuffer_buf(7));
  drc_bufs19121 : INVD4BWP7T port map(I => n_1304, ZN => framebuffer_buf(6));
  drc_bufs19127 : INVD4BWP7T port map(I => n_1310, ZN => framebuffer_buf(5));
  drc_bufs19133 : INVD4BWP7T port map(I => n_1316, ZN => framebuffer_buf(4));
  drc_bufs19139 : INVD4BWP7T port map(I => n_1322, ZN => framebuffer_buf(3));
  drc_bufs19145 : INVD4BWP7T port map(I => n_1328, ZN => framebuffer_buf(2));
  drc_bufs19151 : INVD4BWP7T port map(I => n_1334, ZN => framebuffer_buf(1));
  drc_bufs19157 : INVD4BWP7T port map(I => n_1340, ZN => framebuffer_buf(0));
  drc_bufs19163 : INVD4BWP7T port map(I => n_1346, ZN => calc_buf_out(23));
  drc_bufs19169 : INVD4BWP7T port map(I => n_1352, ZN => calc_buf_out(22));
  drc_bufs19175 : INVD4BWP7T port map(I => n_1358, ZN => calc_buf_out(21));
  drc_bufs19181 : INVD4BWP7T port map(I => n_1364, ZN => calc_buf_out(20));
  drc_bufs19187 : INVD4BWP7T port map(I => n_1370, ZN => calc_buf_out(19));
  drc_bufs19193 : INVD4BWP7T port map(I => n_1376, ZN => calc_buf_out(18));
  drc_bufs19199 : INVD4BWP7T port map(I => n_1382, ZN => calc_buf_out(17));
  drc_bufs19205 : INVD4BWP7T port map(I => n_1388, ZN => calc_buf_out(16));
  drc_bufs19211 : INVD4BWP7T port map(I => n_1394, ZN => calc_buf_out(15));
  drc_bufs19217 : INVD4BWP7T port map(I => n_1400, ZN => calc_buf_out(14));
  drc_bufs19223 : INVD4BWP7T port map(I => n_1406, ZN => calc_buf_out(13));
  drc_bufs19229 : INVD4BWP7T port map(I => n_1412, ZN => calc_buf_out(12));
  drc_bufs19235 : INVD4BWP7T port map(I => n_1418, ZN => calc_buf_out(11));
  drc_bufs19241 : INVD4BWP7T port map(I => n_1424, ZN => calc_buf_out(10));
  drc_bufs19247 : INVD4BWP7T port map(I => n_1430, ZN => calc_buf_out(9));
  drc_bufs19253 : INVD4BWP7T port map(I => n_1436, ZN => calc_buf_out(8));
  drc_bufs19259 : INVD4BWP7T port map(I => n_1442, ZN => calc_buf_out(7));
  drc_bufs19265 : INVD4BWP7T port map(I => n_1448, ZN => calc_buf_out(6));
  drc_bufs19271 : INVD4BWP7T port map(I => n_1454, ZN => calc_buf_out(5));
  drc_bufs19277 : INVD4BWP7T port map(I => n_1460, ZN => calc_buf_out(4));
  drc_bufs19283 : INVD4BWP7T port map(I => n_1466, ZN => calc_buf_out(3));
  drc_bufs19289 : INVD4BWP7T port map(I => n_1472, ZN => calc_buf_out(2));
  drc_bufs19295 : INVD4BWP7T port map(I => n_1478, ZN => calc_buf_out(1));
  counter_reg_3 : DFKCND1BWP7T port map(CP => clk, CN => new_counter(3), D => n_355, Q => counter(3), QN => n_1);
  counter_reg_4 : DFKCND1BWP7T port map(CP => clk, CN => new_counter(4), D => n_355, Q => counter(4), QN => n_13);
  counter_reg_5 : DFKCND1BWP7T port map(CP => clk, CN => new_counter(5), D => n_355, Q => counter(5), QN => n_299);
  counter_reg_2 : DFKCND1BWP7T port map(CP => clk, CN => new_counter(2), D => n_355, Q => counter(2), QN => n_74);
  calc_buf_out_reg_0 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(0), E => n_355, Q => calc_buf_out_0_3514, QN => n_392);
  framebuffer_buf_reg_157 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(157), E => n_347, Q => framebuffer_buf_157_3695, QN => n_398);
  framebuffer_buf_reg_156 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(156), E => n_349, Q => framebuffer_buf_156_3694, QN => n_404);
  framebuffer_buf_reg_155 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(155), E => n_347, Q => framebuffer_buf_155_3693, QN => n_410);
  framebuffer_buf_reg_154 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(154), E => n_349, Q => framebuffer_buf_154_3692, QN => n_416);
  framebuffer_buf_reg_153 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(153), E => n_360, Q => framebuffer_buf_153_3691, QN => n_422);
  framebuffer_buf_reg_152 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(152), E => n_356, Q => framebuffer_buf_152_3690, QN => n_428);
  framebuffer_buf_reg_151 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(151), E => n_347, Q => framebuffer_buf_151_3689, QN => n_434);
  framebuffer_buf_reg_150 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(150), E => n_355, Q => framebuffer_buf_150_3688, QN => n_440);
  framebuffer_buf_reg_149 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(149), E => n_360, Q => framebuffer_buf_149_3687, QN => n_446);
  framebuffer_buf_reg_148 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(148), E => n_356, Q => framebuffer_buf_148_3686, QN => n_452);
  framebuffer_buf_reg_147 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(147), E => n_347, Q => framebuffer_buf_147_3685, QN => n_458);
  framebuffer_buf_reg_146 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(146), E => n_357, Q => framebuffer_buf_146_3684, QN => n_464);
  framebuffer_buf_reg_145 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(145), E => n_357, Q => framebuffer_buf_145_3683, QN => n_470);
  framebuffer_buf_reg_144 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(144), E => n_356, Q => framebuffer_buf_144_3682, QN => n_476);
  framebuffer_buf_reg_143 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(143), E => n_356, Q => framebuffer_buf_143_3681, QN => n_482);
  framebuffer_buf_reg_142 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(142), E => n_355, Q => framebuffer_buf_142_3680, QN => n_488);
  framebuffer_buf_reg_141 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(141), E => n_357, Q => framebuffer_buf_141_3679, QN => n_494);
  framebuffer_buf_reg_140 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(140), E => n_357, Q => framebuffer_buf_140_3678, QN => n_500);
  framebuffer_buf_reg_139 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(139), E => n_357, Q => framebuffer_buf_139_3677, QN => n_506);
  framebuffer_buf_reg_138 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(138), E => n_356, Q => framebuffer_buf_138_3676, QN => n_512);
  framebuffer_buf_reg_137 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(137), E => n_360, Q => framebuffer_buf_137_3675, QN => n_518);
  framebuffer_buf_reg_136 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(136), E => n_356, Q => framebuffer_buf_136_3674, QN => n_524);
  framebuffer_buf_reg_135 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(135), E => n_347, Q => framebuffer_buf_135_3673, QN => n_530);
  framebuffer_buf_reg_134 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(134), E => n_347, Q => framebuffer_buf_134_3672, QN => n_536);
  framebuffer_buf_reg_133 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(133), E => n_347, Q => framebuffer_buf_133_3671, QN => n_542);
  framebuffer_buf_reg_132 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(132), E => n_357, Q => framebuffer_buf_132_3670, QN => n_548);
  framebuffer_buf_reg_131 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(131), E => n_355, Q => framebuffer_buf_131_3669, QN => n_554);
  framebuffer_buf_reg_130 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(130), E => n_356, Q => framebuffer_buf_130_3668, QN => n_560);
  framebuffer_buf_reg_129 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(129), E => n_357, Q => framebuffer_buf_129_3667, QN => n_566);
  framebuffer_buf_reg_128 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(128), E => n_356, Q => framebuffer_buf_128_3666, QN => n_572);
  framebuffer_buf_reg_127 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(127), E => n_349, Q => framebuffer_buf_127_3665, QN => n_578);
  framebuffer_buf_reg_126 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(126), E => n_356, Q => framebuffer_buf_126_3664, QN => n_584);
  framebuffer_buf_reg_125 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(125), E => n_349, Q => framebuffer_buf_125_3663, QN => n_590);
  framebuffer_buf_reg_124 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(124), E => n_349, Q => framebuffer_buf_124_3662, QN => n_596);
  framebuffer_buf_reg_123 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(123), E => n_347, Q => framebuffer_buf_123_3661, QN => n_602);
  framebuffer_buf_reg_122 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(122), E => n_349, Q => framebuffer_buf_122_3660, QN => n_608);
  framebuffer_buf_reg_121 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(121), E => n_347, Q => framebuffer_buf_121_3659, QN => n_614);
  framebuffer_buf_reg_120 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(120), E => n_349, Q => framebuffer_buf_120_3658, QN => n_620);
  framebuffer_buf_reg_119 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(119), E => n_357, Q => framebuffer_buf_119_3657, QN => n_626);
  framebuffer_buf_reg_118 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(118), E => n_357, Q => framebuffer_buf_118_3656, QN => n_632);
  framebuffer_buf_reg_117 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(117), E => n_355, Q => framebuffer_buf_117_3655, QN => n_638);
  framebuffer_buf_reg_116 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(116), E => n_349, Q => framebuffer_buf_116_3654, QN => n_644);
  framebuffer_buf_reg_115 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(115), E => n_356, Q => framebuffer_buf_115_3653, QN => n_650);
  framebuffer_buf_reg_114 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(114), E => n_347, Q => framebuffer_buf_114_3652, QN => n_656);
  framebuffer_buf_reg_113 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(113), E => n_360, Q => framebuffer_buf_113_3651, QN => n_662);
  framebuffer_buf_reg_112 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(112), E => n_356, Q => framebuffer_buf_112_3650, QN => n_668);
  framebuffer_buf_reg_111 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(111), E => n_355, Q => framebuffer_buf_111_3649, QN => n_674);
  framebuffer_buf_reg_110 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(110), E => n_347, Q => framebuffer_buf_110_3648, QN => n_680);
  framebuffer_buf_reg_109 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(109), E => n_360, Q => framebuffer_buf_109_3647, QN => n_686);
  framebuffer_buf_reg_108 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(108), E => n_355, Q => framebuffer_buf_108_3646, QN => n_692);
  framebuffer_buf_reg_107 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(107), E => n_356, Q => framebuffer_buf_107_3645, QN => n_698);
  framebuffer_buf_reg_106 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(106), E => n_355, Q => framebuffer_buf_106_3644, QN => n_704);
  framebuffer_buf_reg_105 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(105), E => n_355, Q => framebuffer_buf_105_3643, QN => n_710);
  framebuffer_buf_reg_104 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(104), E => n_356, Q => framebuffer_buf_104_3642, QN => n_716);
  framebuffer_buf_reg_103 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(103), E => n_355, Q => framebuffer_buf_103_3641, QN => n_722);
  framebuffer_buf_reg_102 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(102), E => n_349, Q => framebuffer_buf_102_3640, QN => n_728);
  framebuffer_buf_reg_101 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(101), E => n_347, Q => framebuffer_buf_101_3639, QN => n_734);
  framebuffer_buf_reg_100 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(100), E => n_349, Q => framebuffer_buf_100_3638, QN => n_740);
  framebuffer_buf_reg_99 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(99), E => n_349, Q => framebuffer_buf_99_3637, QN => n_746);
  framebuffer_buf_reg_98 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(98), E => n_349, Q => framebuffer_buf_98_3636, QN => n_752);
  framebuffer_buf_reg_97 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(97), E => n_356, Q => framebuffer_buf_97_3635, QN => n_758);
  framebuffer_buf_reg_96 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(96), E => n_357, Q => framebuffer_buf_96_3634, QN => n_764);
  framebuffer_buf_reg_95 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(95), E => n_355, Q => framebuffer_buf_95_3633, QN => n_770);
  framebuffer_buf_reg_94 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(94), E => n_349, Q => framebuffer_buf_94_3632, QN => n_776);
  framebuffer_buf_reg_93 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(93), E => n_349, Q => framebuffer_buf_93_3631, QN => n_782);
  framebuffer_buf_reg_92 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(92), E => n_357, Q => framebuffer_buf_92_3630, QN => n_788);
  framebuffer_buf_reg_91 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(91), E => n_349, Q => framebuffer_buf_91_3629, QN => n_794);
  framebuffer_buf_reg_90 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(90), E => n_347, Q => framebuffer_buf_90_3628, QN => n_800);
  framebuffer_buf_reg_89 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(89), E => n_357, Q => framebuffer_buf_89_3627, QN => n_806);
  framebuffer_buf_reg_88 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(88), E => n_347, Q => framebuffer_buf_88_3626, QN => n_812);
  framebuffer_buf_reg_87 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(87), E => n_355, Q => framebuffer_buf_87_3625, QN => n_818);
  framebuffer_buf_reg_86 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(86), E => n_347, Q => framebuffer_buf_86_3624, QN => n_824);
  framebuffer_buf_reg_85 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(85), E => n_347, Q => framebuffer_buf_85_3623, QN => n_830);
  framebuffer_buf_reg_84 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(84), E => n_347, Q => framebuffer_buf_84_3622, QN => n_836);
  framebuffer_buf_reg_83 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(83), E => n_356, Q => framebuffer_buf_83_3621, QN => n_842);
  framebuffer_buf_reg_82 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(82), E => n_356, Q => framebuffer_buf_82_3620, QN => n_848);
  framebuffer_buf_reg_81 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(81), E => n_347, Q => framebuffer_buf_81_3619, QN => n_854);
  framebuffer_buf_reg_80 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(80), E => n_347, Q => framebuffer_buf_80_3618, QN => n_860);
  framebuffer_buf_reg_79 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(79), E => n_355, Q => framebuffer_buf_79_3617, QN => n_866);
  framebuffer_buf_reg_78 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(78), E => n_357, Q => framebuffer_buf_78_3616, QN => n_872);
  framebuffer_buf_reg_77 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(77), E => n_357, Q => framebuffer_buf_77_3615, QN => n_878);
  framebuffer_buf_reg_76 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(76), E => n_355, Q => framebuffer_buf_76_3614, QN => n_884);
  framebuffer_buf_reg_75 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(75), E => n_360, Q => framebuffer_buf_75_3613, QN => n_890);
  framebuffer_buf_reg_74 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(74), E => n_347, Q => framebuffer_buf_74_3612, QN => n_896);
  framebuffer_buf_reg_73 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(73), E => n_356, Q => framebuffer_buf_73_3611, QN => n_902);
  framebuffer_buf_reg_72 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(72), E => n_355, Q => framebuffer_buf_72_3610, QN => n_908);
  framebuffer_buf_reg_71 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(71), E => n_357, Q => framebuffer_buf_71_3609, QN => n_914);
  framebuffer_buf_reg_70 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(70), E => n_356, Q => framebuffer_buf_70_3608, QN => n_920);
  framebuffer_buf_reg_69 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(69), E => n_349, Q => framebuffer_buf_69_3607, QN => n_926);
  framebuffer_buf_reg_68 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(68), E => n_360, Q => framebuffer_buf_68_3606, QN => n_932);
  framebuffer_buf_reg_67 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(67), E => n_360, Q => framebuffer_buf_67_3605, QN => n_938);
  framebuffer_buf_reg_66 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(66), E => n_355, Q => framebuffer_buf_66_3604, QN => n_944);
  framebuffer_buf_reg_65 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(65), E => n_356, Q => framebuffer_buf_65_3603, QN => n_950);
  framebuffer_buf_reg_64 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(64), E => n_360, Q => framebuffer_buf_64_3602, QN => n_956);
  framebuffer_buf_reg_63 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(63), E => n_360, Q => framebuffer_buf_63_3601, QN => n_962);
  framebuffer_buf_reg_62 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(62), E => n_349, Q => framebuffer_buf_62_3600, QN => n_968);
  framebuffer_buf_reg_61 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(61), E => n_360, Q => framebuffer_buf_61_3599, QN => n_974);
  framebuffer_buf_reg_60 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(60), E => n_355, Q => framebuffer_buf_60_3598, QN => n_980);
  framebuffer_buf_reg_59 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(59), E => n_355, Q => framebuffer_buf_59_3597, QN => n_986);
  framebuffer_buf_reg_58 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(58), E => n_360, Q => framebuffer_buf_58_3596, QN => n_992);
  framebuffer_buf_reg_57 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(57), E => n_360, Q => framebuffer_buf_57_3595, QN => n_998);
  framebuffer_buf_reg_56 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(56), E => n_360, Q => framebuffer_buf_56_3594, QN => n_1004);
  framebuffer_buf_reg_55 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(55), E => n_349, Q => framebuffer_buf_55_3593, QN => n_1010);
  framebuffer_buf_reg_54 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(54), E => n_360, Q => framebuffer_buf_54_3592, QN => n_1016);
  framebuffer_buf_reg_53 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(53), E => n_355, Q => framebuffer_buf_53_3591, QN => n_1022);
  framebuffer_buf_reg_52 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(52), E => n_360, Q => framebuffer_buf_52_3590, QN => n_1028);
  framebuffer_buf_reg_51 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(51), E => n_360, Q => framebuffer_buf_51_3589, QN => n_1034);
  framebuffer_buf_reg_50 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(50), E => n_360, Q => framebuffer_buf_50_3588, QN => n_1040);
  framebuffer_buf_reg_49 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(49), E => n_356, Q => framebuffer_buf_49_3587, QN => n_1046);
  framebuffer_buf_reg_48 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(48), E => n_356, Q => framebuffer_buf_48_3586, QN => n_1052);
  framebuffer_buf_reg_47 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(47), E => n_360, Q => framebuffer_buf_47_3585, QN => n_1058);
  framebuffer_buf_reg_46 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(46), E => n_360, Q => framebuffer_buf_46_3584, QN => n_1064);
  framebuffer_buf_reg_45 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(45), E => n_349, Q => framebuffer_buf_45_3583, QN => n_1070);
  framebuffer_buf_reg_44 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(44), E => n_360, Q => framebuffer_buf_44_3582, QN => n_1076);
  framebuffer_buf_reg_43 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(43), E => n_349, Q => framebuffer_buf_43_3581, QN => n_1082);
  framebuffer_buf_reg_42 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(42), E => n_357, Q => framebuffer_buf_42_3580, QN => n_1088);
  framebuffer_buf_reg_41 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(41), E => n_356, Q => framebuffer_buf_41_3579, QN => n_1094);
  framebuffer_buf_reg_40 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(40), E => n_357, Q => framebuffer_buf_40_3578, QN => n_1100);
  framebuffer_buf_reg_39 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(39), E => n_355, Q => framebuffer_buf_39_3577, QN => n_1106);
  framebuffer_buf_reg_38 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(38), E => n_357, Q => framebuffer_buf_38_3576, QN => n_1112);
  framebuffer_buf_reg_37 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(37), E => n_356, Q => framebuffer_buf_37_3575, QN => n_1118);
  framebuffer_buf_reg_36 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(36), E => n_355, Q => framebuffer_buf_36_3574, QN => n_1124);
  framebuffer_buf_reg_35 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(35), E => n_356, Q => framebuffer_buf_35_3573, QN => n_1130);
  framebuffer_buf_reg_34 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(34), E => n_360, Q => framebuffer_buf_34_3572, QN => n_1136);
  framebuffer_buf_reg_33 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(33), E => n_347, Q => framebuffer_buf_33_3571, QN => n_1142);
  framebuffer_buf_reg_32 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(32), E => n_360, Q => framebuffer_buf_32_3570, QN => n_1148);
  framebuffer_buf_reg_31 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(31), E => n_357, Q => framebuffer_buf_31_3569, QN => n_1154);
  framebuffer_buf_reg_30 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(30), E => n_357, Q => framebuffer_buf_30_3568, QN => n_1160);
  framebuffer_buf_reg_29 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(29), E => n_347, Q => framebuffer_buf_29_3567, QN => n_1166);
  framebuffer_buf_reg_28 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(28), E => n_347, Q => framebuffer_buf_28_3566, QN => n_1172);
  framebuffer_buf_reg_27 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(27), E => n_355, Q => framebuffer_buf_27_3565, QN => n_1178);
  framebuffer_buf_reg_26 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(26), E => n_355, Q => framebuffer_buf_26_3564, QN => n_1184);
  framebuffer_buf_reg_25 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(25), E => n_357, Q => framebuffer_buf_25_3563, QN => n_1190);
  framebuffer_buf_reg_24 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(24), E => n_356, Q => framebuffer_buf_24_3562, QN => n_1196);
  framebuffer_buf_reg_23 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(23), E => n_349, Q => framebuffer_buf_23_3561, QN => n_1202);
  framebuffer_buf_reg_22 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(22), E => n_349, Q => framebuffer_buf_22_3560, QN => n_1208);
  framebuffer_buf_reg_21 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(21), E => n_357, Q => framebuffer_buf_21_3559, QN => n_1214);
  framebuffer_buf_reg_20 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(20), E => n_349, Q => framebuffer_buf_20_3558, QN => n_1220);
  framebuffer_buf_reg_19 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(19), E => n_356, Q => framebuffer_buf_19_3557, QN => n_1226);
  framebuffer_buf_reg_18 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(18), E => n_357, Q => framebuffer_buf_18_3556, QN => n_1232);
  framebuffer_buf_reg_17 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(17), E => n_357, Q => framebuffer_buf_17_3555, QN => n_1238);
  framebuffer_buf_reg_16 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(16), E => n_355, Q => framebuffer_buf_16_3554, QN => n_1244);
  framebuffer_buf_reg_15 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(15), E => n_357, Q => framebuffer_buf_15_3553, QN => n_1250);
  framebuffer_buf_reg_14 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(14), E => n_357, Q => framebuffer_buf_14_3552, QN => n_1256);
  framebuffer_buf_reg_13 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(13), E => n_349, Q => framebuffer_buf_13_3551, QN => n_1262);
  framebuffer_buf_reg_12 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(12), E => n_347, Q => framebuffer_buf_12_3550, QN => n_1268);
  framebuffer_buf_reg_11 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(11), E => n_349, Q => framebuffer_buf_11_3549, QN => n_1274);
  framebuffer_buf_reg_10 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(10), E => n_360, Q => framebuffer_buf_10_3548, QN => n_1280);
  framebuffer_buf_reg_9 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(9), E => n_360, Q => framebuffer_buf_9_3547, QN => n_1286);
  framebuffer_buf_reg_8 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(8), E => n_355, Q => framebuffer_buf_8_3546, QN => n_1292);
  framebuffer_buf_reg_7 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(7), E => n_357, Q => framebuffer_buf_7_3545, QN => n_1298);
  framebuffer_buf_reg_6 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(6), E => n_360, Q => framebuffer_buf_6_3544, QN => n_1304);
  framebuffer_buf_reg_5 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(5), E => n_356, Q => framebuffer_buf_5_3543, QN => n_1310);
  framebuffer_buf_reg_4 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(4), E => n_360, Q => framebuffer_buf_4_3542, QN => n_1316);
  framebuffer_buf_reg_3 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(3), E => n_360, Q => framebuffer_buf_3_3541, QN => n_1322);
  framebuffer_buf_reg_2 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(2), E => n_356, Q => framebuffer_buf_2_3540, QN => n_1328);
  framebuffer_buf_reg_1 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(1), E => n_347, Q => framebuffer_buf_1_3539, QN => n_1334);
  framebuffer_buf_reg_0 : EDFD0BWP7T port map(CP => clk, D => new_framebuffer_buf(0), E => n_360, Q => framebuffer_buf_0_3538, QN => n_1340);
  calc_buf_out_reg_23 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(23), E => n_360, Q => calc_buf_out_23_3537, QN => n_1346);
  calc_buf_out_reg_22 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(22), E => n_357, Q => calc_buf_out_22_3536, QN => n_1352);
  calc_buf_out_reg_21 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(21), E => n_349, Q => calc_buf_out_21_3535, QN => n_1358);
  calc_buf_out_reg_20 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(20), E => n_349, Q => calc_buf_out_20_3534, QN => n_1364);
  calc_buf_out_reg_19 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(19), E => n_356, Q => calc_buf_out_19_3533, QN => n_1370);
  calc_buf_out_reg_18 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(18), E => n_356, Q => calc_buf_out_18_3532, QN => n_1376);
  calc_buf_out_reg_17 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(17), E => n_355, Q => calc_buf_out_17_3531, QN => n_1382);
  calc_buf_out_reg_16 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(16), E => n_347, Q => calc_buf_out_16_3530, QN => n_1388);
  calc_buf_out_reg_15 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(15), E => n_357, Q => calc_buf_out_15_3529, QN => n_1394);
  calc_buf_out_reg_14 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(14), E => n_349, Q => calc_buf_out_14_3528, QN => n_1400);
  calc_buf_out_reg_13 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(13), E => n_349, Q => calc_buf_out_13_3527, QN => n_1406);
  calc_buf_out_reg_12 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(12), E => n_360, Q => calc_buf_out_12_3526, QN => n_1412);
  calc_buf_out_reg_11 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(11), E => n_355, Q => calc_buf_out_11_3525, QN => n_1418);
  calc_buf_out_reg_10 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(10), E => n_349, Q => calc_buf_out_10_3524, QN => n_1424);
  calc_buf_out_reg_9 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(9), E => n_360, Q => calc_buf_out_9_3523, QN => n_1430);
  calc_buf_out_reg_8 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(8), E => n_356, Q => calc_buf_out_8_3522, QN => n_1436);
  calc_buf_out_reg_7 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(7), E => n_347, Q => calc_buf_out_7_3521, QN => n_1442);
  calc_buf_out_reg_6 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(6), E => n_357, Q => calc_buf_out_6_3520, QN => n_1448);
  calc_buf_out_reg_5 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(5), E => n_357, Q => calc_buf_out_5_3519, QN => n_1454);
  calc_buf_out_reg_4 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(4), E => n_349, Q => calc_buf_out_4_3518, QN => n_1460);
  calc_buf_out_reg_3 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(3), E => n_356, Q => calc_buf_out_3_3517, QN => n_1466);
  calc_buf_out_reg_2 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(2), E => n_357, Q => calc_buf_out_2_3516, QN => n_1472);
  calc_buf_out_reg_1 : EDFD0BWP7T port map(CP => clk, D => new_calc_buf_out(1), E => n_355, Q => calc_buf_out_1_3515, QN => n_1478);
  g19672 : IND2D1BWP7T port map(A1 => n_302, B1 => counter(6), ZN => n_1482);
  g19673 : IND2D1BWP7T port map(A1 => n_93, B1 => n_59, ZN => n_1483);
  g19674 : IND4D0BWP7T port map(A1 => n_43, B1 => n_33, B2 => n_73, B3 => n_72, ZN => n_1484);

end synthesised;
