configuration memory_synthesised_cfg of memory is
   for synthesised
   end for;
end memory_synthesised_cfg;
