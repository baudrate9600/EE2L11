library IEEE;
use IEEE.std_logic_1164.ALL;

entity gen25mhz is
   port(clk50mhz : in  std_logic;
				clk25mhz : out std_logic);
end gen25mhz;

